module testbench_just_read();

localparam KEY_WIDTH = 32;
localparam DATA_WIDTH = 30;
localparam NUMBER_OF_TABLES = 8;
localparam HASH_TABLE_MAX_SIZE = 11;

reg clk;
reg reset;
reg [2+KEY_WIDTH+DATA_WIDTH-1:0] data_i;
reg ready_i;
reg valid_i;
wire ready_o;
wire valid_o;
wire [2+KEY_WIDTH+DATA_WIDTH-1:0] data_o;

wire [KEY_WIDTH-1:0]                                    logic_matrix [NUMBER_OF_TABLES-1:0][HASH_TABLE_MAX_SIZE-1:0];
wire [NUMBER_OF_TABLES*HASH_TABLE_MAX_SIZE*KEY_WIDTH-1:0]    matrixes_o;

axi_wrapper #(
    .KEY_WIDTH(32),
    .DATA_WIDTH(30),
    .NUMBER_OF_TABLES(8),
    .HASH_TABLE_MAX_SIZE(11),
    .HASH_TABLE_SIZE({256'h0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b}),
    .BUCKET_SIZE(2))
the_table ( 
    .clk(clk),
    .reset(reset),
    .data_i(data_i),
    .ready_i(ready_i),
    .valid_i(valid_i),
    .matrixes_i(matrixes_o),
    .ready_o(ready_o),
    .valid_o(valid_o),
    .data_o(data_o));
    
integer i;    
initial begin
    clk = 0;
    reset = 1;
    #5;
    clk = 1;
    #5;
    clk = 0;
    reset = 0;
    #5;
    for(i = 0; i<100; i = i+1) begin
        clk = ~clk;
        #5;
    end
end

initial begin
    data_i = 0;
    valid_i = 1;
    ready_i = 1;
    data_i = {2'b10, 32'b000000, 30'd0};
    #10;/*
    valid_i = 1;
    data_i = {2'b10, 32'b000000, 30'd1};
    #10;
    data_i = {2'b10, 32'b001000, 30'ha};
    #10;
    data_i = {2'b10, 32'b010000, 30'd3};
    #10;
    data_i = {2'b10, 32'b011000, 30'd4};
    #10;
    data_i = {2'b10, 32'b100000, 30'd5};
    #10;
    data_i = {2'b10, 32'b101000, 30'd6};
    #10;
    data_i = {2'b10, 32'b001010, 30'hb};
    #10;
    data_i = {2'b10, 32'b000100, 30'd7};

    #10;
    data_i = {2'b11, 32'b001000, 30'd0};
    #10;
    data_i = {2'b10, 32'b001110, 30'd2};

    #10;
    data_i = {2'b10, 32'b110000, 30'd8};
    #10;
    data_i = {2'b10, 32'b000010, 30'd9};

    #10;

    data_i = {2'b01, 32'b000010, 30'hff};
    #10;
    data_i = {2'b01, 32'b110000, 30'hff};
    #10;
    data_i = {2'b01, 32'b000100, 30'hff};
    #10;
    data_i = {2'b01, 32'b101000, 30'hff};
    #10;
    data_i = {2'b01, 32'b100000, 30'hff};
    #10;
    data_i = {2'b01, 32'b011000, 30'hff};
    #10;
    data_i = {2'b01, 32'b010000, 30'hff};
    #10;
    data_i = {2'b01, 32'b001110, 30'hff};
    #10;
    data_i = {2'b01, 32'b000000, 30'hff};
    
    #10;*/


    #50;
    $finish;    
end



















localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd11,32'd11,32'd11,32'd11,
                                                             32'd11,32'd11,32'd11,32'd11};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = 
                                                                                    '{'{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001}, 
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001}};

assign logic_matrix = Q_MATRIX;

genvar l,k;
generate
    for (l = 0; l < NUMBER_OF_TABLES; l++) begin
        for (k = 0; k < HASH_TABLE_MAX_SIZE; k++) begin
            assign matrixes_o[(l * HASH_TABLE_MAX_SIZE * KEY_WIDTH) + (k * KEY_WIDTH) +: KEY_WIDTH] = logic_matrix[l][k];
        end
    end
endgenerate













endmodule
