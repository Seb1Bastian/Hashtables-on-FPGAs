module matrix_generator #(parameter NUMBER_OF_TABLES = 4,
                          parameter HASH_ADR_WIDTH   = 5,
                          parameter KEY_WIDTH = 6)(
    output  wire  [NUMBER_OF_TABLES*HASH_ADR_WIDTH*KEY_WIDTH-1:0]  matrixes_o
); 

wire[KEY_WIDTH-1:0] logic_matrix[NUMBER_OF_TABLES-1:0][HASH_ADR_WIDTH-1:0];

localparam [KEY_WIDTH-1:0] Q_MATRIX[31:0][16:0] = 
              '{'{64'b0010101011111011101010110100000111010111011111011001110100010100,
                  64'b0010100011010010100111101011110011011011001000101110001111100101,
                  64'b0001001101011110011111101010000110011101101011111010110000001100,
                  64'b1011101001011000101010110000011100111001111011110110001000111100,
                  64'b0010011111101000011010101100001010100000100001101101000000000011,
                  64'b0110111011101010111100110011010001011101101001100100101101100011,
                  64'b1000001100000101111101111001011010001010010101111010000110101101,
                  64'b0001000011001110100101111010010001010101011001010111110010111001,
                  64'b0000101100011001101010010010101011111000100111001010110111010101,
                  64'b1011111100101101011100000111110011111011101001010111010101101000,
                  64'b1011110101101010001100100101100111011000101011010000010001101101,
                  64'b0101001101000000001111101010000101101000101111001010111000011110,
                  64'b0110101011100000011010000011000011000011011110111100111100011000,
                  64'b0111000010011000001101010110001011100111101110001001000111000100,
                  64'b1010001110110001010101000110001000011000100100111011000101100110,
                  64'b0111110001100010010101001000000010111000111010000100010000001001,
                  64'b1011011111011110010100010010111111000011111001000101001101001110},

                //30
                '{64'b1111011010111110010110100000111110010010000000101101101100101100,
                  64'b0010110010101111110000111100101111100110110010100011110111101011,
                  64'b0010000001110000010100000011111100000000011100111001100101110110,
                  64'b0011111001001110110001011111010010100101011001101101000011011110,
                  64'b1111000100111110011000101111011101010000101111010010011110100000,
                  64'b1010000010100111001101011110111001110001010100011101011011010111,
                  64'b1110011011000010111010011101100011011111111001110011011101010111,
                  64'b1101111101000101001111011110110101111001010010000001001010111100,
                  64'b0000110100001010101000011101001011011010101101101001110100010110,
                  64'b0101001000101011010100110011001001000001010011000000001000110001,
                  64'b0001100100100110110001111010010010111001110111001001011110000010,
                  64'b1110110010011110010111000000101101101110111011010010010010100100,
                  64'b0011011100001000010011000100011100110111111101100111100010001100,
                  64'b1100000010101010111111000100101011110101101010001011010110111000,
                  64'b1000010110000101011010011010000101011011000001000011100111011011,
                  64'b0110000110001100000100000101011100011111110111000000001011111111,
                  64'b0101000000100110101101100000111000000100100011001100000000011101},

                  //29
                '{64'b0111110100101101111100001101001010100001010010110101001100011000,
                  64'b1101100110101001111100111111011111000011010001001101010001010100,
                  64'b0100111100000111010001100111101101001100011110101101011011110011,
                  64'b0111001110010101100101100101011001111110000100100001000101111011,
                  64'b0000000111011111101000011001000100111010010110101001111001100111,
                  64'b1011111001010100100010010011010110101111000111110010001000111000,
                  64'b1100010011100010000010010111111100111011010111101010110101011111,
                  64'b1110000110011010110000111001111100000110100110011100011010101010,
                  64'b0011100111000010011101011010110011001010100011100010001010001010,
                  64'b1111100111111111010101100111000010110010011010010000110110101001,
                  64'b0100010011111001000000101101100110000110111110111011011001001101,
                  64'b0101010001001010111100011100101111001000000111101001011101011101,
                  64'b0100110011000000110011011110001111100001011101110110100010110010,
                  64'b0000110101011100111111111100011111101111110000010011011110110001,
                  64'b1110010101111110010010011101000101000110000001101011001001000001,
                  64'b1001001101111011100011001011010001100011101100010100001000011101,
                  64'b0001001010010101011010000011011110001110101000010001100001100110},

                  //28
                '{64'b1101101100010011000000100100010111101101010000110101000010111110,
                  64'b0100011000100011010101100100000011100000000100110011110010011000,
                  64'b0010011011010100100110001100110101010101010001000111100010110001,
                  64'b1110110000100000010001010000100100101011110111110100001111001001,
                  64'b1111001011000011101101111110100100110100011100000000011101010011,
                  64'b1100010111010011100110000110100010101100100010011100010011110110,
                  64'b0110011110011110100000111110000111100110000001111000000000001100,
                  64'b0000110001000110111111010110001111101000111100111000100111111001,
                  64'b1010000101100011101101111110011110001111101101000101100011011100,
                  64'b0101011111010110100010011111011001000010111011101111111110111001,
                  64'b0100001111001110111111000001100101001000101111011111010110011101,
                  64'b0000001100111101110101000111000010000111111111010111100110000101,
                  64'b1010010101010110111010011011110101010000000001110011110101110010,
                  64'b0101000010111100100001110111010110100100100011110111011111010111,
                  64'b1011010010011011000001001011110000001111010000100110101100011111,
                  64'b0001111100111100111111101010100011010001010001010100101001000101,
                  64'b0010011110100110010000111011010000011100100111100110111010101010},

                  //27
                '{64'b0010101001001001000001000101011001011100010111000101101011010110,
                  64'b0001011111001111110101100100001001000100010000101100001001111001,
                  64'b0100111011010111101100100010000100100101000110111001110101000000,
                  64'b0010111110010011001111000000111001000111111101100000000001011010,
                  64'b0011101101000011110101101111001111001001101001000101000011101101,
                  64'b1101001000101011011111000101010100101111011001001011111010000011,
                  64'b0111101000100000110001000110001001001000001110000111000111010011,
                  64'b0100101010010011011101110001001110110101101111100011110101011011,
                  64'b0011010000110001011000000010111100011110000100100101000101000010,
                  64'b1000011110110011011001100011000101011111111100101011110011111101,
                  64'b1011111100111100000000010000001010101110011011101001110010001101,
                  64'b0100101000010001000011001001001011010010000010011110010000000011,
                  64'b0010100010100010010100011111010110011001100000000011000100111101,
                  64'b1101100010110111110000110000010110001110111000100110100000101110,
                  64'b0110110111010001110100001100100110000011111011100101110101111101,
                  64'b1001000010011011101111100010010111100001001000010110100001000100,
                  64'b1011110011000001001110111000110110011101101111000110111011000000},

                  //26
                '{64'b0111001010100001000100110101110001000010011010111011000011111001,
                  64'b1111011001111001010101101001110101000000001001001101111101111011,
                  64'b0100011010111111011101110010101000010100000011101101110000000000,
                  64'b0001010000110111100000111110101101010010100111010011010110100011,
                  64'b1011010000010100110101010010110101100111011110010101100100011111,
                  64'b0001101000001000000111111010100010000110111001000001110011110001,
                  64'b0011001110101101001100011011011110001100011111101010111001010100,
                  64'b0000000111110111001110010101010100101010110011100111010001101010,
                  64'b0011111111111110010000010100000010000101011010100111111110011100,
                  64'b1110100010000001101111111000110110110000111010010100101110111010,
                  64'b1101000101100101101011000110100100110101000000011110111000011100,
                  64'b0100000001010101001100000100000111010001000110011011000000111110,
                  64'b0010100100110001001111000010111001011101011100101101010001010111,
                  64'b0011101000101111011101011000111101111101110101000110101111100011,
                  64'b1100111001001010011000010001000101010111010111011110011000100011,
                  64'b1110000110111001000001101110011001001000101010100001100000101011,
                  64'b0011011000010000110011111100011010110110111100001101110011010111},

                  //25
                '{64'b0001101101011001100011101010000000000110101011110010110111000000,
                  64'b1100011011011011101101111010111001011110101110111010101000011111,
                  64'b1000111001101111000010010110010001101100011010000010100011100000,
                  64'b1110010000011101100000101011100000101001110100000100111001101100,
                  64'b1010010010001010010111010011000100100110010110010000000010111010,
                  64'b0000010010101010000011110110000000001011100011001110011101010000,
                  64'b0111111101101110101011110001011100110000100010011000010001111101,
                  64'b0010001011000000111101110000101110110100101011001100001010111101,
                  64'b1000000001010001011000001111110000010101010111101100101101000111,
                  64'b0111000011010110011010001110001111111100010011001000111111001100,
                  64'b0111101101110100001100010100000011000110110001101010111001110010,
                  64'b0011111101110110001001011001001010111000000000101101011111100111,
                  64'b0101111001000001010111111100110111111010100100010110011100101010,
                  64'b1000000011111110000011010000010110000100100100110101100110010010,
                  64'b1110100001011010110010111000010101111110000111011000110101001001,
                  64'b1110001000000000010101100010001101100111011101110110110010111101,
                  64'b1100110100000100000010000100110100110011111110001000111000101001},

                  //24
                '{64'b1010110010111100011000011000001001010110101011000000010111101100,
                  64'b0000010001010001110011100000110101010001011110011000110001010000,
                  64'b1110100111110001110011110001110110100011011100001010101111110101,
                  64'b1101001011111111100001010000011011111110111010100010100010111101,
                  64'b1001000110111111111110101100011010011000111001111100100011011110,
                  64'b0010111001011110100000101100011101100010111010000111000110010110,
                  64'b1100011111101001010010110101100100011000001011010010011100001010,
                  64'b0111001001000001100011100100110001001101110011000110000101000001,
                  64'b0010111011001011100100100100110011100000100110110011010111011001,
                  64'b0101110101000101011111001010001100001111111000101000010101111010,
                  64'b0011111011101011000110110110000000111001110100110010111111101110,
                  64'b0110011001010101001111110010111000110101011000001101011100111110,
                  64'b0011000000001110101110111110111111011010011110111001101000101000,
                  64'b0001001110100111100100010000011111111110011010110110010101111011,
                  64'b0000110110110100011000100111101100100000100110111010010111010110,
                  64'b0000111110100111110001001100000110110110011111111111100100101100,
                  64'b1111010001110101001011111001000111000111010011000111101001001001},


                  //23
                '{64'b1010001011000100010100110110110000111000010000101001100100010111,
                  64'b0100001001011001010101100100111011110111001001001000010000001001,
                  64'b1010000000110011000111001000111101100100000010101111011101111000,
                  64'b0110100000010101011011000101010100011011011100110001010000101011,
                  64'b0001010011111110010110001100111011110111000100101101101001000101,
                  64'b0001100101110101110100100110011011100010010000001111000100100101,
                  64'b0111001001111010101110100010111011101100011100101100111010011100,
                  64'b1110010101110110011000111001001000100000110011001000000000110001,
                  64'b0110010110000100110111000001000110011001100111100110001000100100,
                  64'b1111101011010111001011010001010110000010000101110010001011001011,
                  64'b1010011111001000011001110000101111101110010101101000110110010110,
                  64'b1010101000100110100000110010100101001001011010011111001100000100,
                  64'b0101100001110111110110010011110100111001000000111011100010100011,
                  64'b0011110110101111000000010000000010110000110110011000001010100100,
                  64'b0111010111011011111101000110000111111011000100110111000100000000,
                  64'b1111010110111111110100101010010111101001001010101110111010101110,
                  64'b1110000000111010001011110100010101100010011110011000001100111000},

                  //22
                '{64'b1000100011101101000001100110111011000010100110101001000110100101,
                  64'b0001111011101010001101010111111101110111100010011111010101100001,
                  64'b1000101011110011111100100001000101011001101011101011001110000101,
                  64'b1100111111101100111111011100000010000100111000000010000110101111,
                  64'b0010001010010001100110010101011000000011010000100001101010010101,
                  64'b0111110100000001110011010101101111000111110101101011001010001100,
                  64'b0000001111011001011011100011101111101111110101011101110101110100,
                  64'b1101010000010111101111000100111100100101110101100111000001110110,
                  64'b0000100010110000010011101110100010010011011100111110011100001000,
                  64'b1101101110110100101110111101101000101010001111101110010000100001,
                  64'b0011100110101010011110111110011101000011111100010101100001001011,
                  64'b0010000111111101001010111100000000011100111111101011011011100100,
                  64'b1110100011010010011010100111111010110010000011110110111111101110,
                  64'b0111000110111011010000101010011001111101110110000001010110001000,
                  64'b1110110100011000111110000111010100100000011111011100110110001100,
                  64'b1011001001011101101000000010111101000011000011100010010001001011,
                  64'b1101011110111110010101010011111000000100101100010001110110011000},

                  //21
                '{64'b1010100111101000101110010000100100011011100011001001010101000010,
                  64'b0011110100001010000111110110001100110001001000010101101010110010,
                  64'b1010100111110001001011001001000110101010101110111000101101111011,
                  64'b1101101010100111011110110101100101110110100100101000001111101001,
                  64'b1100000100100001111110110101010011100101110101101101010111101000,
                  64'b0111100010101111100110011101100001101110011101000010110101000111,
                  64'b0000101011000000110111111000100111100001101100011110100100000001,
                  64'b1001000111101001010101000011111010011000001011000101101000111011,
                  64'b1000011001110101011010100100011000100100100000100110100111001100,
                  64'b0010000010100111111001010101110101010111010010111010110110101011,
                  64'b1001100010110011101111101010110101111110100100111000001101100101,
                  64'b1110001011110110001011101010110111011001001110110110110010110100,
                  64'b0010011111101011111111110000110101001001101000110100100101011001,
                  64'b1011010110000110100000001110110101100111010000000111001000000011,
                  64'b0011001001110100010111001110000100000100101011001100011010010111,
                  64'b1010110110101010101000101100100000001001101011100010110101110110,
                  64'b1010111110100101011000100010101001000111100000100110101000101101},

                  //20
                '{64'b1110001001001001100111111100011110111011111111010010001100100000,
                  64'b0100000001011101111100000001000000111100010111101000001000011000,
                  64'b1101000011011100101011100110011000110010011100010001100000010101,
                  64'b1100011010000010101001011100011111110000101000001000110101011011,
                  64'b0000010111101101101110111000000000010110011010101010100001000111,
                  64'b0111001100101101100101001100000010100000100100100011101010111011,
                  64'b0100110100101101010000100110011100011100011110011110110011100111,
                  64'b0010000111111010101011000001010100110000011110000011000111110111,
                  64'b0000110000101010001111111001001010100000111011001110101100110010,
                  64'b1101011001111011000111001011110001100001100111100000110001001011,
                  64'b0001000010010010101011110111001100100011101000011101000101000101,
                  64'b0010101000010100010000010101100101001011111001101110111101011010,
                  64'b1001010001001000101000000110101111110111000100111011011000000001,
                  64'b1100010000000100001011001000101011101010111001010010110100110101,
                  64'b1101001100010000111110100101010110011110011001100111111101001110,
                  64'b0111110001110110010111011101010001111101010000011101000000100110,
                  64'b1110110011110111111000011101000111010101011000011111110100111010},

                  //19
                '{64'b1111100010111101110010100110000100010011000100100100010110100110,
                  64'b1110011010110100111100110110000111010100011110011001101110010010,
                  64'b1000101110100111101100001001000100010001111011011111110010001110,
                  64'b0100101100111110000111001000011001100100100100000101001010110010,
                  64'b0011111000011001001100010101111101100100110011111110010100111101,
                  64'b0010110010110111100001011101011000100111110100100000110000111110,
                  64'b1011000111101011001000000110111010110111111101011110011101010001,
                  64'b1011001001101010000101111010101001010110000011101111100111000010,
                  64'b1010101000001101000001000110010010001000100011111000111100110100,
                  64'b0010110110100110000101100100101010110010011101110010010100010010,
                  64'b0010001011101001111100001010001010110011010001011010000011101001,
                  64'b0100110001100101010111110011101111101011010010010111101111111010,
                  64'b1001110001100010000101111111110111000110010010010000111101110000,
                  64'b1010011111110011111001111011101101010011000010101010011000111111,
                  64'b1011000100110110010010000001010011100110001111111100110110001011,
                  64'b1110011001100011000111000010010010010001001000001010010010000000,
                  64'b1011101011101101101101110011111010000111110100010111010101100110},


                  //18
                '{64'b0000110001100000001111010100100110101110100100101101111000110110,
                  64'b1111011001100100000110000001011101111110011101111000100001111001,
                  64'b0100011110010101110010110101010100011110110010100100111000001100,
                  64'b1011010101111111110000001011100111111111110010100110001111110010,
                  64'b1100111100000110001011001100010010010100110100100001000010011011,
                  64'b1101001110110000100000111010010110100101100101010011000111110000,
                  64'b1001100001011010100011111000010101010010111011011101101000010001,
                  64'b1111111110101001010001100111100111100100000100110001001001010100,
                  64'b0001011000110100011110010100011010011101110100011000011110010100,
                  64'b1100100011110011010110100011001100010000000011101101111110000100,
                  64'b0100001011110001001110001000000110100111101001001110111011100000,
                  64'b1100111011111010011110000101100100010011100010011000101101101010,
                  64'b1000000111010101100001011011010011000111110101101110011001010100,
                  64'b0000110111100000001001110000010011101101110100101110010000011011,
                  64'b0111110110100001000100000101111101100111111111010110101010010000,
                  64'b0111011000010000011010010111010000010011110110000001101110010011,
                  64'b0110011111111000101001111101110111011100101001111010001111100011},

                //17
                '{64'b1010010010100011100110001110000101011100101111100110111000100001,
                  64'b1011001010110101000110111100010000010011110001101011110111100100,
                  64'b0101110111111100110111011000111010001111100101001111101101111010,
                  64'b1000010011100011000110101000011100000011010011110011101011001000,
                  64'b0101000011100010010101010001011010101011001110111010110101111101,
                  64'b1111010000110000010101110100011110001010100010010001101111000101,
                  64'b1000000000000000110010001111101000100110011000001110001100000010,
                  64'b0010101110101110110111000100001101110001111001000011001101001101,
                  64'b1011010110110111011001100010011100001101101111011000010011011110,
                  64'b1000011000110010011100000000101100001111000101010001010011111010,
                  64'b0000100101100011000101011110010101011111010111101100000100111010,
                  64'b0011001100000000010001100110100100101010011101000011111100001111,
                  64'b0000111100100011010010111110110001001001101111010011101011110010,
                  64'b1001011000101010001101001011011001101100101010010100110111111001,
                  64'b1100001000011001100100101110010111110010100111000000000101111110,
                  64'b0001001101101001100111110001110011010000011111000001010000111010,
                  64'b0100001101100111001000101000101101000000101000011000011010100000},


                  //16
                '{64'b1001111010101001001100010001000111110001110110110100101100000011,
                  64'b1101111011100010010100011000100110111111010100100010011111010000,
                  64'b0010100100001011001111100010111111010011111011111000010100000110,
                  64'b1110000010110000101000001101010000001101001110011011000010011110,
                  64'b0010111100001101100100110101011101110000010000100100111011101111,
                  64'b0011100010101001101010011100000100001010001111011110110011111010,
                  64'b1001011001011010011000001010011000101101110100011000111011100111,
                  64'b0010100011010110100001110100010111001100010100011011000101011100,
                  64'b0110111001010011101001110100111110000111101101110111101010111110,
                  64'b0111001110010011011101000100100011111101110101111010100111100000,
                  64'b0111110001110011110100010111111100001011110010011000101010000111,
                  64'b0000000111000010010001100100111000101000000101011111010110001100,
                  64'b1000000000000010101000111110100100000001101000010001000100001000,
                  64'b1101100001100011100110100010101111011000001011001101011101101110,
                  64'b0011100010011100111001101101110000110101101010001001101101100000,
                  64'b0111001110011001100001010010110011101001011110110111101101011111,
                  64'b1101010010101101100001011010101001111111011110011100001111011011},

                //15
                '{64'b0000011010111111110110110011011010011001101110000100110000001110,
                  64'b1111110110010101011100011111101001110111000110100010001010111011,
                  64'b0011000010010001010110111111000000110101011010110100000010011000,
                  64'b1011000001010110010110001001110111111011011111000110010001000001,
                  64'b0100001000111000101101001000011011000001110001110000000111011000,
                  64'b0011110100111100111000010101001001011111100010001010001100001000,
                  64'b1101001101000110100111000011111000111111111010010011000111110100,
                  64'b0001001011001001110101010111010011111010010001001010100001000111,
                  64'b1111001001110000011010010101010010101110101011001001001001011010,
                  64'b1110000110010111000010001010000010010010100010110111101010101111,
                  64'b1010110100011100010010110000111111000000111001010010001100001011,
                  64'b1100011100100000010101000101011000111011111100001100000100001000,
                  64'b1001111011010100100001110110001011001101011011100010001110011011,
                  64'b1101100110101011100001000011100001001111001010001000011111101100,
                  64'b1010101111001101000000100111100010000111001110010000001101100101,
                  64'b1110101001001111111011001110001000101110010110111010010011110101,
                  64'b0010101001100101000001100110000100001001110010110111000110101000},


                  //14
                '{64'b0111101010001010110110111110101011110101000111110010010001000011,
                  64'b1000011111110000100010100001110011101001100100101101011110000000,
                  64'b0101100101001011100100100101011011100011100001111110010010100000,
                  64'b0010111110110101111000101000011100011110111110010010110011001111,
                  64'b1001011101011001111110100100010010001100111010010100110000111000,
                  64'b0001110100000110000000011000000011011000011001110100001100011000,
                  64'b0000011010001000111100011111011100111001111110111011100011000001,
                  64'b0010001011110000000111111001100001111110110111010111110000011010,
                  64'b0100100100010100100101011011010111001000101001010100010011001011,
                  64'b1001111010011111111001111111101001010011000110100110101101110011,
                  64'b0011000100011100001001011110000001010001010010001111010011100110,
                  64'b0001100101101001111100010001111011110011001000001100110101110000,
                  64'b0001101010100100011001100110100110100011101110011101110011001111,
                  64'b1001101100110101100001010111110010000110110010101010100010110111,
                  64'b1100110101001010101111000111111001010001001111000100001100010010,
                  64'b0110101001000011101010011010010101101111101111010101000011001100,
                  64'b0000010110001001000111100011011011010101000101011000101110100100},

                //13
                '{64'b0010001110100110010001111111101001000011010011011101000010001100,
                  64'b1110011111101101110100000011111111110111101110101000100111111000,
                  64'b0010101101110110001111111100110100101110101001110000100011001011,
                  64'b0101000000110100101010100100010001010001011000110010010010100111,
                  64'b0111100011001001010101100010101001000010001001111011100110011010,
                  64'b0011101111101011011100100110100100101101110110111000101101101011,
                  64'b0100100011010001010000000001100111110001111110100011111010100010,
                  64'b1101010111111001101010111000101101001110100011110110001100001100,
                  64'b1001011111010100101100111001100110101101000110001001000010001101,
                  64'b1100111110011101010000110110010010100110110101100001100110001000,
                  64'b1011101100100010100001011101010110000001110100010000010011001000,
                  64'b1001001011011100111100010111101111010110010101010011010111111101,
                  64'b1001100101101010011000110010001110010010000101111001000110101101,
                  64'b0111000000001110001110111101101000000010110110001101111000110010,
                  64'b0101011010011000101100001101000010110001110000100110110101100110,
                  64'b0000111011100110001001110001001100010110111100101111100011001111,
                  64'b0010010100101110110111000000111110010011011101000111100101001101},


                  //12
                '{64'b1110110010101011001011111111100010111000001001011001111110101010,
                  64'b1100111100111010001010010101111010111110010001111011110000001100,
                  64'b0010110101110010110111111101010111110101001011001010001100010000,
                  64'b0111000001010011100111010011111000101000110000001011011101011011,
                  64'b0010110001001111000010100010011100011110100001101000001111110100,
                  64'b1000101100100001000110001110001111111011110101010100100010111110,
                  64'b0010010101101101000001110000001001101001101000000100100111101000,
                  64'b0000011110101011000111000111010100001101001000001011111000100000,
                  64'b0101101100100001010110110101000011010001100100000101000010010100,
                  64'b0010101110010101001100001011011011110111100111011000100001010011,
                  64'b1110111110001101111100111010011010100011010111000001001000010100,
                  64'b0010001010001110101010001000100011110111110101000110100010000100,
                  64'b0011001111101110000001100001101011110111010101011010100010000011,
                  64'b0010011000001000110001111100110011111000111000100101111001011100,
                  64'b0111111000111101010101100011110001100010000010111001010000101011,
                  64'b1110001000001111110011111011000100100101001111111011011100101101,
                  64'b1101110001010001111111000000111010110011010100011100010011101001},

              //11
                '{64'b1000010111111001000001001100011111101101100111010000111111010011,
                  64'b1101000110000111101100000110101110100101001010001000111010100101,
                  64'b1110111111111001000101010010100011001010101101011100111100000101,
                  64'b1111010000001101111111010100010111010111010100101011000000001101,
                  64'b1010000011000111101101110010100101111001111111110000110101110000,
                  64'b1100000001101000100111010111001110000010111010010010110101111001,
                  64'b1010100011100101001111110010000001100101110100101111101101110001,
                  64'b0000100101100100011110100010000100000111110110011000001001000100,
                  64'b0101011101111101001111100001101110101010001011001001100011000101,
                  64'b1010101101011011001110011011011101111111000101010110111000100001,
                  64'b1101000101000011110010100110000000111111000011001000111101011100,
                  64'b1111001111011010011000110111101000100011101101000100100100111000,
                  64'b0011000111100011010000010111011010010000111001001110001011000010,
                  64'b0110011001001010011010001111000000000111111001100110100011011101,
                  64'b1101110100000100110000110011110001001101010000010111100101011011,
                  64'b1101010110111110010101101010010101111010011110010001110100011010,
                  64'b0000111011100011001011010000000011000011101100110011010001111001},

                  //10
                '{64'b0100101011110010000101010000100111100100011001011011111000110001,
                  64'b1011010111001111110000110010101001001101100001011110110000011010,
                  64'b0000010100100000011101011011100100011010110001000101100110011010,
                  64'b0100100011001111011010001011110000111101110001010011010101000001,
                  64'b1001111111110010000001101001100100000010001111110001011011010010,
                  64'b1001111001111011001001000000001110001011011000110100001111111100,
                  64'b0111100110000001011001110001110010101100011001011111110001011110,
                  64'b0001001110101001010011001010100110010110010110000111101101010100,
                  64'b1101100111000111000001101010001011010110111010101111011011000110,
                  64'b0110111010010010000101101100001111010111001110011101001110000110,
                  64'b1100010111010000101001110111110101111101101000100111101011101110,
                  64'b0010101110010100111011101110111111001110100011010101100010111000,
                  64'b0100011111101001111111011100101111111111000010111110100111101010,
                  64'b1101000001001000010101000011001111001101100000010101001010101001,
                  64'b1001111000110000110010101100000100111100101101100001110010110111,
                  64'b0100010000000101111010111110000010010111100100001011000000111000,
                  64'b0001011001110100100011110001001001000001010111101010010101011111},

              //9
                '{64'b1001111001100000101100101000011011100100111011100111010100001111,
                  64'b1010000000001000100100101111111010110000101000100001100101111011,
                  64'b0110110011100100000010011001100010001001010010110010010110100001,
                  64'b0111011011101010000100111110110111111110001001010001111110100001,
                  64'b0101010110110100001011100011101001110001111110100000011001100001,
                  64'b1010101100001101001011111010110010101100011101001110010101011110,
                  64'b0100110111010111000101100111111000100110001000011000100011001101,
                  64'b0011100000000000010001011101010000001110010001100100000010001011,
                  64'b0100110101010001011110011001000110011101111011110011011010111111,
                  64'b0101101011101111101100010010010110000101100110000101001101111101,
                  64'b1001010111010111110111001011111011011100000010100011011001110111,
                  64'b0000101000011011111110110011010010000000110000100101100111000100,
                  64'b1010011011000011100101000101110001110101110101001101101000001111,
                  64'b0101110001101000110011110110011010000000011001010101101000110111,
                  64'b1001001011101011101000010001010010010111110100111100110011011111,
                  64'b0100111001010001111000001100011100111110011101110011011101010110,
                  64'b1001010110000011111111101010111000010010001000001000001001001011},

                  //8
                '{64'b0000000100001001101011000010010101111000111011101010011010110111,
                  64'b0010000111011101110011111110100111110000110110010011110000100111,
                  64'b0100010010101100101110100001101101011110100111001000000010001100,
                  64'b1100011111100100101110000000000110001100000101010111111001101001,
                  64'b1101110110101110110010011010011011001001001000011110100110010010,
                  64'b0101111010011111111100100001011101010111001011011011011010100100,
                  64'b0000010100000000111011100110100010100110110110000011111101001010,
                  64'b0100011000001101010101100000001010001101110000100101001111101011,
                  64'b0010110101100001101010011001000110001111011111110010010100111101,
                  64'b1101111001011001100111101001111101011111001100101000110110000010,
                  64'b1010111100110110111101101100010010001111111010101101100011100011,
                  64'b0110000101000010010110001000010110001111000100011011011110100100,
                  64'b1000001111100001101001111101101001001011001111000110011001101101,
                  64'b0001011000101011110011101101110000110100100100100100101001001010,
                  64'b0111010111110000001100110100011101000110101111000010110011111001,
                  64'b1101011001110011101110011000001111001101000001001000011101010100,
                  64'b0101000100110111010100001011110001101011100100100100001001101100},

              //7
                '{64'b0101101110110001100011010011010011010110101101011100010110010111,
                  64'b0110010110111111010000001000111101111000001011111101100001111110,
                  64'b1101011010110001011001111111001000001100111000011111101111011000,
                  64'b1101100000000101110001000010111000001101010110011001011110101000,
                  64'b1001111111011011010001011010100010000101010011000000011101001100,
                  64'b0000011101110010000001011101100101110010111101011011101011100011,
                  64'b1001011001001101111011111101010101101001111101000000110101010110,
                  64'b0100001010011001001011000100110111110001111100110101101110010000,
                  64'b0111010111011110101000111011011010101010000010111000001101101010,
                  64'b1101010100001010011111111011100001100010000101111111001011011000,
                  64'b1111011111000011001110110101110010000000011001001111100000000000,
                  64'b0011011100001110000110010101011101001001110000101110000001101111,
                  64'b1100100110101111000100000001100100001010001101011101011011011011,
                  64'b1010100110110000001111100101010000101010101001111011010110100111,
                  64'b0010001110100011111110011110110101010010100101001000110111001011,
                  64'b0111100001000010101111111100101111010010010010011110010001101001,
                  64'b0000110010110010110100111101011110100111101011110010011010011100},

                  //6
                '{64'b0000001100001000000011111101010101010000010000111111110110101001,
                  64'b1000101101110110100110110001101000111101010011010010100100001001,
                  64'b1011010001011010000011111000110010011010110110011110010101001111,
                  64'b0011110000100100101100111110011000010100010001011010001001111000,
                  64'b1111111100011111111000011110010001011101100011010111010000110000,
                  64'b1011010011010011011010010000011111101001110011100000110101101010,
                  64'b0100001110001101011011000110010000001011000000011011000110010011,
                  64'b1110010001100101111100100111000001110100110101111101000100100011,
                  64'b1010001011100011001100000000110000111011001110101110010111001111,
                  64'b0001101111010100100101110111011000111000010101110111111011101101,
                  64'b1110011110110111001011011101111001111111010010110000101101011110,
                  64'b1000010001111011111011001110101011001100011010111100101101001001,
                  64'b0100101101100011000000001110000010101011110100001100100010100001,
                  64'b1011010110010110010011111101111110001101100000011000010011110000,
                  64'b0000010100001111001111110000100100011011110011011111011100010000,
                  64'b1001101110011100001101100101100100011000110011100011111100111111,
                  64'b1011001111010111000001111011001101111010101011111111100001101001},

              //5
                '{64'b0010101110011110110011111011001101100010011110110111010101111000,
                  64'b1110101111011001111011011111101011000010011010100011110101010110,
                  64'b1100100001001110000111110110111011100100000110110000001001000111,
                  64'b0011011100010011111011111111111111110111010011011111011100100100,
                  64'b0101010001111101001001110111110111110111110101010011100000101101,
                  64'b0111111001100110011111111010101100110101001010011111000011000010,
                  64'b1010010110010010011001101000111011111011111010110011011111110100,
                  64'b1110111010000000001001010000100011001111110000010111001011011001,
                  64'b0000001001101101101000000110000011111100100101010001010111000001,
                  64'b1111101111011101000011001010010100110011011101100111000110110110,
                  64'b0101000111011010010010100010011010001101001011011000110100100000,
                  64'b1000010011000111101001001100100010101011010000100010010111010011,
                  64'b1110001111001100011100111101101101111110101010001100011101011010,
                  64'b1111111110101000000100100011111101010000000100000100010101101001,
                  64'b0100001110110101001011100101110010111101111110110000000110101001,
                  64'b0000010000000100110000110011100010000011001001010111101001010101,
                  64'b1111111001111001100111100110110100001011101110010101000010010100},

                  //4
                '{64'b0110001110111000110001000011000110110110010101101011111100000001,
                  64'b1001010111010011001101111001111101111000000101000010110100000111,
                  64'b0011100100000111101111010100001110101110001011010011010011001100,
                  64'b0111111101010001010101000001001001101100110111001110100010100011,
                  64'b0100011110010111111101100010100100101101001111000110100001101111,
                  64'b1000111101000101011111001001001010111110110010111111011101011101,
                  64'b1001000100101100100110000110100101000000000011010001010000111001,
                  64'b0101100000011101100010101011010011101110011011010101100010010110,
                  64'b0110010111011110110000100101011101100001101100100110011100100001,
                  64'b0111110001001010100111101011001000110111111100110001010001110111,
                  64'b1111000101111010011111001010000010001110010101010011010100010001,
                  64'b1011011101111100011101001110110011111010110010011111111010010101,
                  64'b0011001100111111111111010111100110011100100110101010100010001101,
                  64'b0111111110011111110110000001000000110010110111101000101001111000,
                  64'b0110011010111110001100101011000111011001100011111110000100011011,
                  64'b0000001000010010010011110010111000110001101101110001110000110000,
                  64'b0001001011000001000111111101001010100101010000100011011001000101},

              //3
                '{64'b0100010101010001000010101100111011101100000001110001110101010000,
                  64'b0001010111111010011100001111100110011001111111101010001101011001,
                  64'b1001111001111011100110101010011100100110010010111000011101001111,
                  64'b0111001110100001010110011101101010001001111110101000011101101011,
                  64'b0111110101100111010001101110001010110100111101000101010000101010,
                  64'b0100101110011100101101000100101001100111000111000100110110100110,
                  64'b1111010110101110011001011100101100101001001100101110100110011010,
                  64'b1010111101010111010001110101011101111000110111000111110101000101,
                  64'b1011001010100011101001111110100101101100101000010100101011110011,
                  64'b0001001001010001000100011101110110100001010101001001001010110101,
                  64'b0001011011111000110010101111010110100000101011011001110110100000,
                  64'b0110010001010011111111101010100100001100111100101110001010101111,
                  64'b1110101111101011110110000101011101011101011000000011000111010100,
                  64'b0011000001110101000001101110111001100111100100010011101000001100,
                  64'b1101110001001011101010110011011110100001001011110010110011101010,
                  64'b0011111011000101001101110110101010101011100010111101100100010100,
                  64'b1110011111101001111000110000001100100111110000100011000000011111},

                  //2
                '{64'b0110111011010110101010010110110111101110100101100111010110111100,
                  64'b1101010111000111111010110111001011011101001111000100101110101011,
                  64'b0111011100010111010101011110100000001101101101110001011010110001,
                  64'b1000001100110001000110110101101000001101010000111011111110111110,
                  64'b1110000111100110101110100100101001110110110111010101100001110110,
                  64'b1100101011011001110101110100001000110100000110000000100110000000,
                  64'b1111100001000000100111010010111110100110100111011111011011100100,
                  64'b0010001000111101001111111110110010000111000000111011000100011001,
                  64'b1011000000001101010100101101111111010111000110101011011110110110,
                  64'b1000001100101000010011001011111101100001000000001101111000101100,
                  64'b1001101111100000111001010011110000101011100110000101000110000110,
                  64'b1010101110111001011010101100110100101100111001011000101011100111,
                  64'b0111001000111110110100101010010010110101111100001111000000111101,
                  64'b0010010001001000110111111111100110010100101010110010101101001001,
                  64'b0101101110100100101000010100001001010110001010010111101110011000,
                  64'b0110001110010000110110110011101100011110101111100000111011101011,
                  64'b0101111010100010100101110110111111110001100001001101101011101001},

                  //1
                '{64'b0101110100010010000100100000100010111011001010100110011011100100,
                  64'b0010000110000011010100000011001010100100000100101101001011101110,
                  64'b0010110100011100100001111010011101110011011100011011101110100111,
                  64'b1000110111111111101001110001001101100000011111010100001001010010,
                  64'b1011010001100101111010101011001001000010001111001100000101110010,
                  64'b0010010010001000101000110111000111111111011111011011100000000100,
                  64'b1011000100000111011001000110110001111110111101111101110000000100,
                  64'b1110100111010011110110000111111001110100010011111101100010000001,
                  64'b1011101000110000101101100001001110101111000001000010110010100110,
                  64'b1001001011011001010000100000111100011100001110110100011001110011,
                  64'b0011001000110110011010101101001110011111100101011110100111100010,
                  64'b1111101110000011011000001110101000011101111100001110100010010101,
                  64'b1010001111010101010001011001010010101001111110110100100000011101,
                  64'b0000110011000111000000000010001100010100110000001101101010001010,
                  64'b0101001101000010001111110001000001110000100011011010101000000000,
                  64'b1111101100010001110100110110001001101010111000000001111111011000,
                  64'b1000011110110001000101101000111110000011000111000001111011111111},

              //0
                '{64'b1101110111011011000001101011110001110100001001000001111101100101,
                  64'b0000101111010101101000011101000010001110000111101011001111110011,
                  64'b1100101001001111111111000111101111110001111000010100000001101100,
                  64'b1000000001101001000011010101011000000111010101001001001011000100,
                  64'b0101111010101001101000011110010011101111100110111000010111011011,
                  64'b1011111100011101101000101000011111111010110011100111001000110000,
                  64'b1101110000111110100010001110100101000101011101101101010001111000,
                  64'b0111000010010010111001110110000111101010010010001000101010000001,
                  64'b1011100011011001111000111111010110100100111011100011000000010100,
                  64'b0110110001111000010100100011010111111110001001000001100101100110,
                  64'b1000000100001101010110000101101000011110100111011000110000100011,
                  64'b1100111000011110111100001101110010101011000001101001010001110110,
                  64'b1110111101011011001100000111011111001100001110100011100101011111,
                  64'b1111110011011011010111101101111100111111011001100101000010101110,
                  64'b0110101100111110010111011000101001100010010101011001010000010111,
                  64'b0001110110010101011100110100110100101100100000000010010111000010,
                  64'b0101101000101101101111000111010110010101010001010101010001100000}};


                  
                           
                                                                                      
genvar i,j,l;
generate
    for (i = 0; i < NUMBER_OF_TABLES; i++) begin
        for (j = 0; j < HASH_ADR_WIDTH; j++) begin
            for (l = 0; l < KEY_WIDTH; l++) begin
                assign logic_matrix[i][j][l] = Q_MATRIX[i][j][l];
            end
        end
    end
endgenerate

generate
    for (i = 0; i < NUMBER_OF_TABLES; i++) begin
        for (j = 0; j < HASH_ADR_WIDTH; j++) begin
            assign matrixes_o[(i * HASH_ADR_WIDTH * KEY_WIDTH) + (j * KEY_WIDTH) +: KEY_WIDTH] = logic_matrix[i][j];
        end
    end
endgenerate

endmodule