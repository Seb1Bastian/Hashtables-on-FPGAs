module matrix_generator #(parameter NUMBER_OF_TABLES = 4,
                          parameter HASH_ADR_WIDTH   = 5,
                          parameter KEY_WIDTH = 6)(
    output  wire  [NUMBER_OF_TABLES*HASH_ADR_WIDTH*KEY_WIDTH-1:0]  matrixes_o
); 

wire[KEY_WIDTH-1:0] logic_matrix[NUMBER_OF_TABLES-1:0][HASH_ADR_WIDTH-1:0];

localparam [150-1:0] Q_MATRIX[7:0][16:0] = 
              '{'{150'b010010100011010010101011010001001001100101100110010101100000111010011111110111101101101100011001100101110110111000111001011000110000111000111110100100,
                  150'b100100000011100000101011100111010111111010010001001011001011111010101001011111010010101111000010101010101100010011110001111000010101101111111100010101,
                  150'b011001101010010001110011010111100101001100000101011001001010010101001110011000010001001101001000111011101110100000000010110000001100011110110001001011,
                  150'b010001011000001111110001001111001010101100111010111110011100011010110011110111101100000000011100000011010010100001000101011011001110111111101011111010,
                  150'b100010101111111110000011100100100001001000010010101010010101001000001000000001011010111010111010010000001101111100100001000101001001011011000101011011,
                  150'b001100110110100011000011111000110011011101100100011011010000111001010000110101010111111010000111001111011110010011010000000010100111100011111010010101,
                  150'b001011001011101101011110110110100111100011011011110010011010111001011110000010010001100010010110100011110010101101101010100010010001010100011111101111,
                  150'b000011001110011000110011110111110000101100100111010111011011000111101101010101100001011001000001101100100101010100101011110111100100101110000000100001,
                  150'b101110110010010000100101001010100100111100110101100010011111110101000011111111011110110101110000100111010010011000011011001001010100011010000001101111,
                  150'b110111001101000110101000100010001110001101001101101110111000001000111010011010110000001011101101010111100101011001001111100010100110111111110101111110,
                  150'b111101001101101001110010010101111100010001100001100001110111010000010110100101111001010100101100110011010100011001000011000001010110110000000000000101,
                  150'b001100010111100001110011110000010111011001110110000101011001100100010110110000111001110010111110111001011000000110110010111010001100001011011011011001,
                  150'b011101010101110001001111111011110001000011111111000101101111100000010011100111101001101110101010111100010100111000011010010000011101010001001011111000,
                  150'b001111010110101010010100011011110001111111011110010100110000101110001000000011101110001000110101000101111100101000100010100010000111101101010000100010,
                  150'b000001010111000101010001010101111111011111001110100110011001100011110100000110011001110000010001100110100010100100001101001100001010111000101010110011,
                  150'b010000011101111011010110100000110000111110001010010000110001001101010011000100110010010100001100010001010110101100110011110010101000011001110111000101,
                  150'b011111100011110110110001100101110011100001111000110100101010010100100101011111110101110000011010011111000111001101110001110010111000010001010011000000},

                //6
                '{150'b011110011001111101100011000100100000101001100000100001010101110010100000101111100100111111100011110111000010100111110111101110100000000011111000010011,
                  150'b100111000001011100101110101011001110011100010010010101011000001111000011110110111100111101101110001110010101100110110110111101110110011010111001101000,
                  150'b100110011100111111010010010111010110001101111011100110001111001010000101100010001101110110010010110001110111101100001011010000011100110110000011111010,
                  150'b111110101011110101001010001000010001001001000101111011100101010000100001110010101101111111111110000010101101010010101101001110111011000111111001111000,
                  150'b100010001100010011110011111011010010110001110001100000000111101011000001011001100000100001111000011001110010110000111111011111011000010110111101100010,
                  150'b111100110111101001111111100000010111000000001001110010010111100101001001100110111100010111000010011110001100011110010010101111101011110111111011011101,
                  150'b011001000100110111101110000011011001110001111011010100100011101100000001110011100011110101000111110000011010010011010101010101000000011001001101011011,
                  150'b100111010100001000001100010011010000010000111100111000111010110101100011110100110101010110111010100110011110110010010111110110010001111000001101111001,
                  150'b110100010111100011000100111100001000011110110101010111111100101000011000101010000111011111011011011101101111001111001000010110100001100100101011001001,
                  150'b111110010100111000011000110111001111111101100001010011110110011000001011101100100111001101000110010101010001110100110011111110101110000101001000001100,
                  150'b010110100100111100000111101011001000110100111000110100111101101010111000001101110101011011000101011011010011100010110111010111101010100001011011000111,
                  150'b000100011011010101001101001110010100110101100010000010001101001111100011111011011100000011110100110011001011100010111010100010011110111010001011011100,
                  150'b111110110101011101000001010011101111010011011011100101101111000011111111000101110001100011011101011100011100011011101001101000100000110100100100001101,
                  150'b001001001000000000000110111101111010101011101010000110000111101111010101100000001100111110100110010000000110001111010001001011010111110100100001111100,
                  150'b000111101111101000000111110110010100010000101101111011000011000000011101000111101010010111111101001011011011001011001110100010110100000100011101101110,
                  150'b101010010010010111101000110010101111001100010111010001110110000000001111011000101100100011101001001110101010101001101001101011100000110110100000100010,
                  150'b110110010110100100011000010100010000001011000001100101101000100000010111000000101000100111000000110011111011001001100110101010001110100100001110101100},

                  //5
                '{150'b001110001000011100110011110001000011101011100101100010000000011101100001001101011100100011110010110100001100000100001010110010011111001111110010111001,
                  150'b011001010111101000101010100010011110000010011100100010001010010000101111110111110100011010001111101001101100011011011100110000010010110010011010100111,
                  150'b100111111001010101000100000100101000011001001111001000101011101100011010100011000011110111000100111001101101000111110000001101101000111111110101001000,
                  150'b110000011100100000001011010111011111000001001011101111011010110011100111000100000101010000111011111111000110001111011010000011111000100101000101011101,
                  150'b110011010101111000000001101010101110100111010110100010101111101100011011001011011000011101100110010011101011100000110110111111001011010100100000011100,
                  150'b101100001111101101111100100010101010101000001101001111000100111000011100000111011101011100110000101001001110111111001100010110101000011010110101101101,
                  150'b011000010001011110000100000111111011101011010010100001010110101101010010111010110000000101111101111101100001111101010010110001110010010000111000000111,
                  150'b101100010011000110011111100011110101010011101010110101110011111001100000111111101110010100011111110111111010110100111001001111000010001011110111011000,
                  150'b111011010001011010111100001010001101011110100001000101011110001010011111100010110111111001001000000000011110111011110001101000101111000000001000001010,
                  150'b100100011110011011100100001101000101010100000000000001110011111001101001011110000111111000110111011001110010011001100111001100101011100100110101101110,
                  150'b110100100000100010100001101000011000101010110010010010000010010110101011111000110011111000001100011110100111101010010000011110001100010101001101110111,
                  150'b000000100111011100001111000111011110100010101001100110010011101000100000011111010011010010000101000001000101110110101000111001011000001001100001110100,
                  150'b100000011111010110000011110000000010101011000100000101100100101111100011000101011001110100111101110100000110100000001011011111100011011111010001000100,
                  150'b100100101010100000111011101001100000001110011011110110101110111010110101101010010001001011011000110010001100011011010101110011100110011011000110011010,
                  150'b001001010101111101100001101000111101111101000011101100010111010110000100011011111011010011011101001111100110010101111100001010100110100100101000000111,
                  150'b111001011001100010101101111001011111101101000100010100100010101110101011001011100000000011100000101100001110011011001000110110000001000011110110001111,
                  150'b100110011001110111010101011001011100011111001101100011010111010011011001010011001011100001101111011010101100000000100111101000110100111000001011101011},

                  //4
                '{150'b010001000110010101101110011100001010101100011010110011011001000000011110111101011110100110001111100101010100110001011011100010010110001011001011001110,
                  150'b101001010110010000101000001001111101011111000101111111011111101110011000011100110111000101010011110110001100100001010010010101111110101110110101100011,
                  150'b010100010000110011010111101001000110100011101011001110000101010001110111100110101101101101011001011111010100001111111001001110011100011011010110110010,
                  150'b001111110001110001001010000000011010101111101000001101010000001001010010111011101110000101111110100000000101111011101101110101011000110001101100100101,
                  150'b010110101111110011001001001100110111010110111010100110110100101110011001101010110101010101110000000110111110110111011001110001010001000101001110000100,
                  150'b000110111100110001110111010000111101000110000010001010100111011011010100110010100001010100001011101101001101010111010111001101100101100011000110100000,
                  150'b111110001001101011110001101000110110011000011010111110010110000101001011011110100101101001010000100110101001110111000101100101010010000101110011111000,
                  150'b101101010111010111101110110100101011110010110101100100001001100010001011111111111100000000100000111001101111111010011010011101000111110101111000011111,
                  150'b010101011111010010110110101101111011010111110110110001010100111100011111011110111011000110001110011100011000100001100010100010101001110101110111110001,
                  150'b110101001000010111101100000000000001011100011010011001011000011010101011110100110101100100011011001011001110010011100110100101110110101111111000010000,
                  150'b100001010001100110010011001111011000100011111101000000001110011111100101001000010010011111011000110010010011110110010101010000000100100101100100010101,
                  150'b010110000100110011101100111000100101000010010000111110010100110110101101001101010011111111101011110100110000001111101001001101101011000101101010110100,
                  150'b101011111100101001000011001100011011011010110100010110101100010011100101110001100000001100001000111101011100011011100010001000111101001100001110111000,
                  150'b001100111010000011101010110001100100001011101111010000101011100010100111000111010000100101010010100001001001000111100011001111001010011111101011101001,
                  150'b001011011100101000000101111100101101000010001010010110111110000100100111100101001100111110101101101000111010000101111000001101111010011110011001100101,
                  150'b111111101000001010011001001010000110101001001001100011110011101000000110101000110101001110010000000111010110101111001101011110011100000100001101000011,
                  150'b101000010110000010101101111000100001000110101000101001010000110111001011000010000100111000100111001100100110011101110100110001110110011010000100001001},

                  //3
                '{150'b001101111010100000010110010001011001001100010110111110110011000100110111011001100110100010010111010100001011011011111101001011100011010001011110100001,
                  150'b011111000010000011010101011111111010101100111011111101110111101110110010100100011011110100101001010110111110110010110100001100001110111100000000110111,
                  150'b010000110010011000111110110111100010010111110000111111011010110010111111011111101000101100011011111101110100110101101100010110010110010011001100011110,
                  150'b011101100110010000100011010011100110101100000101000100001101110011011000100001111110111100011001001100111101010110111001010110101000011110111001010101,
                  150'b001001101110010101000011000111110101111001011011111001110000110000001011111000100001111011101111101100001000011000111011101111110100100001100111000000,
                  150'b100011001001011110011110010010110100110000111101010111111110101001001010101001100001111110010010110010010111000010111001001001111010010010001011000100,
                  150'b000010110000111000010100010001010001100000010110100000001011000000011010110011101110101100001000010100101000100110000100000000101010110000100100000000,
                  150'b011001101000100101001101010100011001001101001101101000000010011110111011011101101000111101111111010000000100101101010110110100011010100101010011011000,
                  150'b010100000011100011011101000000100001110101101001101100000011111100001110111010110001001111011101110111010010011101111111101000100100000011110000110111,
                  150'b100011011101010011000110100111100010111111011001000110000011011110101001100011000101100010011000111010101011110101100000011110100001111010011111001001,
                  150'b110010111101010011001101100110110101111001100101011101000101111011000010111011100101000110000011000011010100010101111000111000011100011010111010000011,
                  150'b001100101111110111010101000110011100011110110010101101011011101011101100001001011101001000111110100010010010111010010011100010000100110001010100110001,
                  150'b001111010001001001100101001100110010001101011110100101110101110111110110001111110001000110101001010101110011010111110101011001000110010000111001011000,
                  150'b101110000100011111011011000011000111101000000101001011011000010000011110010001011111000111100110100010011111111011100001100001010000011001100001111111,
                  150'b101101111011000011100011101001010011100111001111010100111011010101101110010010100000101110000101011101001000101000010110101000100111010101101011111011,
                  150'b010000100011110100111010001011110011000100010001100110111101000001110010110100110111110101000111100001001110011010101100110010010000100111010001001110,
                  150'b110101000111011111111000010111001011111110011110111100011111011010000100011110110001100111011111101110010001000111110111001010100011111111010101101111},

                  //2
                '{150'b011001011001111001111110111100111100100110010100001111100001101101110001110001010111110010100101010001011011111011010110001000110010001101001000010010,
                  150'b011110100000011000011100010000111101101110001011101111110110010110110111001111001001111000001100011010011101110101100100011001111110110001100110000001,
                  150'b100011100001101011110011011000111010110010001010100101101001011100101110000000001011010010100000001001001110000100100110100101111000010111111001101010,
                  150'b000100111101011011001111110001001111100100111100001101101101101100011100011100110011101010100100100110101011100010000010101000101001100100110001110111,
                  150'b010010001000000011101101101111010010011011110101101001100001111101010010110111111001010011111100010111001110111011011011001000010001101011101011000101,
                  150'b101010100110100100010011110111111000101101011110110101110011001010111000001101110100111011100111011000010010110111001111111000110011110001110110111110,
                  150'b111000110000110111011101100101010000111010011010100111101111010001110111011000010111111001010011001101101000010111011011010000100011101110011110101010,
                  150'b010001000010011100011010000101011011000111101101111011010011110010101110000110011011110100001101000001000110011101001110010001011111000001001101011111,
                  150'b111010000111010011000010010000000100011000000011111011011001010000011000111110100000011110010100110001000011000001010100101011011000010111010110101101,
                  150'b010101010100101011010001101010010000010000001001110101111010010010101001100000111010110010000111101110110110111100000000111011010011110000100100010100,
                  150'b011000111111111011100111000101011011101000101111001001100101100010110010110001111011100000000011110011010111110110000110000110101100010010011001000100,
                  150'b011101000011010111101101001010001000100010110110100000010010100001001110001101010100110111010001111010000000011110110000100011010000001001001010111101,
                  150'b101101001011101100100111110001010011000001110110001001101011010001001000001001011100001110111010000111110100001110011001110000011000110100000000010000,
                  150'b100000010011100011010100010011011110100111011111001111010110011100110110110101111001000001000101111001011001100101111000111011011111101001101100111000,
                  150'b011001100111001100101110110100110001011001110111011010001000010101111100101100011000111011111100010010101010011011101111010111110110000111010001111111,
                  150'b110011001100011011010100010000111000100111010110011000110110110100011001001001011101101100111101010011000010001000010001101000110101000001110111000110,
                  150'b100110110110011101111001001111000010000000010011111010101000000011111101110100101111010001110101011101110101011000110110010111101110001000010101111110},

                  //1
                '{150'b000011000101110111111000101100101111010110001101010011101011110110001010100101101110110111000000011101011001100100110000111100010010110010101000001011,
                  150'b101101101010001101100101110000001000001010011111111110000011110001001010001010011001001110101110101011000010011111110101011101100111010000100010011100,
                  150'b001001001011111000100110010111110101000110100101001001101011011101110000000110110011100110001100010100111010110101100100101110100101101110001111111001,
                  150'b110010001110101101110110001100011000000101010001101010111101100110101000101100101101110010101110001100011010011100101110011011011011110111011100110111,
                  150'b000111111111001110000100101000100110000001111110010001011010010000001010101100110011101111101011010011000011111110000111100000110000100110001000110000,
                  150'b010100110000001010011101101001110111110100010111100100110011000001110100011010110011000000011010110001100011110010001000001111100010101010110011000100,
                  150'b111011111111110001000111110011100011011110001100001111000001011011011110101000011111111001101001000000100001010011100000001000101110011001111011000111,
                  150'b001111110101001100000111001100000111010111000011010111101010100001100010011110111010111101001011101100010010011101100100111100001110000100111110101110,
                  150'b111000000110001100000101111011110001110111111110101010010110000001101111110101101111110001001011100101111101111100111001010101100001010001001110011000,
                  150'b011000101111010111101100111011110101000110000101011101000110010001111111001111000011101110010100100011101010010010001011111011011000011010011001100001,
                  150'b000100011111001001100101100111100010011011011101111000110110011111100100000111110010010100000011100011001000000111101011100010010111100000101010010100,
                  150'b101010111000001001110101111111101011000100100111101110011110101110001010100100110101010011110100101110000110010111000100000100101001100110101110110011,
                  150'b101011111101100001110001100100001000010101100001110111010000100101100111000001111111101001111110011110101101010110100011010111110100100000100100100111,
                  150'b101010010100100011111101111001100001000000001011100101000001010011100111001110100010111011111110010011001000011110010001100100111100101010100000100111,
                  150'b011101101001100111101000011111111101001010100110000101101111000000001110100101101100101110011101001000110011110111000100111101110010001100111011101011,
                  150'b101001101101010000000111111001110100111011010011111001000001010111110101000010001101110001111100101110110111111111100100000001110011100111011010111100,
                  150'b010111010010000101011011111111010101011000101001101101010101111110100111011101001000110010110000101001101110110001001101010100100001010001110111100000},

                  //0
                '{150'b100001000000100111001101111101010100001110010100001101100001110011000111111010011110011011110001010101111101110110110001101010001110000011000011111101,
                  150'b000100111111011111011010100100010111110110011010000110001000101111001001011101010000011101111110101111001001110010101010101000010011111011101111110010,
                  150'b100111111100110110100110011011101011100100111000110011010000010010110101110001101011111001110111011101101010010000000110000001101010000010000011000100,
                  150'b100001111100011101101010101011001011110111110010011110101101011111100001000010000110000010000000110000011010001100000110011111101001001010101011100010,
                  150'b111010000110111010101000111101101010110101011110110110011011001100011101110101110010011011111101110011110110010101011001100111010011011110001010110111,
                  150'b000010111011101000000010010000000111001000101101000010011100101111101111010000011011011110100100111100100101011010111010000011001100100100010101111010,
                  150'b100101100101111001110010011101101100101100100000110011111110010110100000100100010011111000001110101110110110011000100011000100101001000111100001000010,
                  150'b010001010101111110100110110111010101010111101100000100100111001110000111110101001010010110010001101011001010010101010111011111011111101000011001110000,
                  150'b111000110001000011111010110111100111011000111111110100011100100010011001100011000101011100000110000011010001101000101001110111100001100011001110101101,
                  150'b010010000000010101001011010011110001101001101101110010111011110010110111001111101000010101111001011111011000001001111111001000110111010011101110100111,
                  150'b101010001010101011001100110000001110101101111011111001110110001111010011111001011111100001110011101011001001101100011011011101100001101100101001001101,
                  150'b011000100001010101000010111101100111001010000101010001001010010010101000000000000011011011010001110001111110101110011110110011001000101011111010110011,
                  150'b011000000000011110011110001001011011110110110100100110010111011111011110100010100011100111011110000000010011001101000100111011010001111011100011000101,
                  150'b101100000111100100011111011001011011010001001100000000000100000101110101010000110001000010000000111010000101010101111011101011110110001101011111110101,
                  150'b100111110100111011110100011100011100111110001100101111010110101001011100011100000011101000101010001001011101101000011101011101011010100110111000001110,
                  150'b101110111011110100100001100110111111111010001001001110001010011001010101000010100001010011100111111101001110010000110000111110011110000100001011010100,
                  150'b001001111101000111000001111000101011001000010100001011001001000100011000001001110110001101110100111011000101111101111011011110111110010010011101110111}};



                  
                           
                                                                                      
genvar i,j,l;
generate
    for (i = 0; i < NUMBER_OF_TABLES; i++) begin
        for (j = 0; j < HASH_ADR_WIDTH; j++) begin
            for (l = 0; l < KEY_WIDTH; l++) begin
                assign logic_matrix[i][j][l] = Q_MATRIX[i][j][l];
            end
        end
    end
endgenerate

generate
    for (i = 0; i < NUMBER_OF_TABLES; i++) begin
        for (j = 0; j < HASH_ADR_WIDTH; j++) begin
            assign matrixes_o[(i * HASH_ADR_WIDTH * KEY_WIDTH) + (j * KEY_WIDTH) +: KEY_WIDTH] = logic_matrix[i][j];
        end
    end
endgenerate

endmodule