key: 15, hash:10, tables: 10
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = '{'{15'b001001100011100,
                                                                                        15'b000000000100001,
                                                                                        15'b000000100011101,
                                                                                        15'b100010111010001,
                                                                                        15'b010000011110100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100010011000,
                                                                                        15'b100011100100110,
                                                                                        15'b011001000101000,
                                                                                        15'b111110001001010},
                                                                                    '{15'b010001011001001,
                                                                                        15'b001000000100000,
                                                                                        15'b001000010100101,
                                                                                        15'b011100010001000,
                                                                                        15'b100011110001111,
                                                                                        15'b001000101000100,
                                                                                        15'b000000000011000,
                                                                                        15'b011111000010000,
                                                                                        15'b000001000100101,
                                                                                        15'b000110000101101}, 
                                                                                    '{15'b000110100000110,
                                                                                        15'b101100110000100,
                                                                                        15'b010001001000111,
                                                                                        15'b001110010010100,
                                                                                        15'b101010010000100,
                                                                                        15'b000101101011001,
                                                                                        15'b001011000010010,
                                                                                        15'b110010100010010,
                                                                                        15'b001000100010110,
                                                                                        15'b110001100010000},

                                                                                    '{15'b001001000011100,
                                                                                        15'b101100000100001,
                                                                                        15'b011000001011101,
                                                                                        15'b010010101010001,
                                                                                        15'b010110011010100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100011011000,
                                                                                        15'b100010001101110,
                                                                                        15'b111001000101000,
                                                                                        15'b110010101011010},
                                                                                    '{15'b010001011001011,
                                                                                        15'b001000000111000,
                                                                                        15'b001000010000101,
                                                                                        15'b011100010101000,
                                                                                        15'b111000110001111,
                                                                                        15'b001001001000100,
                                                                                        15'b010001100011000,
                                                                                        15'b011011000000111,
                                                                                        15'b011001010000110,
                                                                                        15'b100100110111001}, 
                                                                                    '{15'b011001100111110,
                                                                                        15'b110110100011010,
                                                                                        15'b001010101000000,
                                                                                        15'b100001101011100,
                                                                                        15'b011111111001000,
                                                                                        15'b110011101110101,
                                                                                        15'b101010110001001,
                                                                                        15'b010000010111011,
                                                                                        15'b000110100110010,
                                                                                        15'b100101011011101},
                                                                                    '{15'b101010001011100,
                                                                                        15'b010110101101000,
                                                                                        15'b111010010000101,
                                                                                        15'b110000111111011,
                                                                                        15'b101100110111000,
                                                                                        15'b110001001010111,
                                                                                        15'b101100110000001,
                                                                                        15'b101001110110010,
                                                                                        15'b010101010111100,
                                                                                        15'b000101011011010},
                                                                                    '{15'b011001000000100,
                                                                                        15'b101100001010000,
                                                                                        15'b000000110101100,
                                                                                        15'b101111110100100,
                                                                                        15'b010011100111000,
                                                                                        15'b001100000001010,
                                                                                        15'b000111101110110,
                                                                                        15'b101010010001011,
                                                                                        15'b000101010110101,
                                                                                        15'b001100011001111}, 
                                                                                    '{15'b110111111011111,
                                                                                        15'b100100111110001,
                                                                                        15'b001011111110100,
                                                                                        15'b110100001010110,
                                                                                        15'b010110011110010,
                                                                                        15'b010001001110100,
                                                                                        15'b100110001011101,
                                                                                        15'b010111111111001,
                                                                                        15'b101000001100001,
                                                                                        15'b110011010111010},
                                                                                    '{15'b101010100101001,
                                                                                        15'b101011111101011,
                                                                                        15'b000011011010100,
                                                                                        15'b110011000101011,
                                                                                        15'b111011000111011,
                                                                                        15'b000001101000100,
                                                                                        15'b111000011100000,
                                                                                        15'b110011010010111,
                                                                                        15'b100000111110111,
                                                                                        15'b101011111010100}};


key: 15, hash:13, tables: 10
localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = '{'{15'b001001100011100,
                                                                                        15'b000000000100001,
                                                                                        15'b000000100011101,
                                                                                        15'b100010111010001,
                                                                                        15'b010000011110100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100010011000,
                                                                                        15'b010011101111010,
                                                                                        15'b100001111000101,
                                                                                        15'b101101111001001,
                                                                                        15'b100011100100110,
                                                                                        15'b011001000101000,
                                                                                        15'b111110001001010},
                                                                                    '{15'b010001011001001,
                                                                                        15'b001000000100000,
                                                                                        15'b001000010100101,
                                                                                        15'b011100010001000,
                                                                                        15'b011100000101100,
                                                                                        15'b001001110100101,
                                                                                        15'b101010010001000,
                                                                                        15'b100011110001111,
                                                                                        15'b001000101000100,
                                                                                        15'b000000000011000,
                                                                                        15'b011111000010000,
                                                                                        15'b000001000100101,
                                                                                        15'b000110000101101}, 
                                                                                    '{15'b000110100000110,
                                                                                        15'b101100110000100,
                                                                                        15'b010001001000111,
                                                                                        15'b001110010010100,
                                                                                        15'b101010010000100,
                                                                                        15'b000101101011001,
                                                                                        15'b001011000010010,
                                                                                        15'b110010100010010,
                                                                                        15'b001000100010110,
                                                                                        15'b001011001110010,
                                                                                        15'b110110101110010,
                                                                                        15'b001011100000110,
                                                                                        15'b110001100010000},

                                                                                    '{15'b001001000011100,
                                                                                        15'b101100000100001,
                                                                                        15'b011000001011101,
                                                                                        15'b010010101010001,
                                                                                        15'b101111000100001,
                                                                                        15'b011001101011101,
                                                                                        15'b110010101010001,
                                                                                        15'b010110011010100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100011011000,
                                                                                        15'b100010001101110,
                                                                                        15'b111001000101000,
                                                                                        15'b110010101011010},
                                                                                    '{15'b010001011001011,
                                                                                        15'b001000000111000,
                                                                                        15'b001000010000101,
                                                                                        15'b011100010101000,
                                                                                        15'b111000111001111,
                                                                                        15'b010110110101000,
                                                                                        15'b111000111010111,
                                                                                        15'b001001001000100,
                                                                                        15'b001001001000100,
                                                                                        15'b010001100011000,
                                                                                        15'b011011000000111,
                                                                                        15'b011001010000110,
                                                                                        15'b100100110111001}, 
                                                                                    '{15'b011001100111110,
                                                                                        15'b110110100011010,
                                                                                        15'b001010101000000,
                                                                                        15'b100001101011100,
                                                                                        15'b011111111001000,
                                                                                        15'b110011101110101,
                                                                                        15'b101010110001001,
                                                                                        15'b101011101110101,
                                                                                        15'b101010110110001,
                                                                                        15'b010011010110011,
                                                                                        15'b010000010111011,
                                                                                        15'b000110100110010,
                                                                                        15'b100101011011101},
                                                                                    '{15'b101010001011100,
                                                                                        15'b010110101101000,
                                                                                        15'b101101110101001,
                                                                                        15'b110101001010110,
                                                                                        15'b101000110011011,
                                                                                        15'b111010010000101,
                                                                                        15'b110000111111011,
                                                                                        15'b101100110111000,
                                                                                        15'b110001001010111,
                                                                                        15'b101100110000001,
                                                                                        15'b101001110110010,
                                                                                        15'b010101010111100,
                                                                                        15'b000101011011010},
                                                                                    '{15'b011001000000100,
                                                                                        15'b101100001010000,
                                                                                        15'b000000110101100,
                                                                                        15'b101111110100100,
                                                                                        15'b010011100111000,
                                                                                        15'b110011110110001,
                                                                                        15'b101101010001010,
                                                                                        15'b100110101110110,
                                                                                        15'b001100000001010,
                                                                                        15'b000111101110110,
                                                                                        15'b101010010001011,
                                                                                        15'b000101010110101,
                                                                                        15'b001100011001111}, 
                                                                                    '{15'b110111111011111,
                                                                                        15'b100100111110001,
                                                                                        15'b110110010110010,
                                                                                        15'b011001001100101,
                                                                                        15'b100101001011101,
                                                                                        15'b001011111110100,
                                                                                        15'b110100001010110,
                                                                                        15'b010110011110010,
                                                                                        15'b010001001110100,
                                                                                        15'b100110001011101,
                                                                                        15'b010111111111001,
                                                                                        15'b101000001100001,
                                                                                        15'b110011010111010},
                                                                                    '{15'b101010100101001,
                                                                                        15'b101011111101011,
                                                                                        15'b000011011010100,
                                                                                        15'b110011000101011,
                                                                                        15'b111011000111011,
                                                                                        15'b101011011100000,
                                                                                        15'b110111010010111,
                                                                                        15'b100100100110111,
                                                                                        15'b000001101000100,
                                                                                        15'b111000011100000,
                                                                                        15'b110011010010111,
                                                                                        15'b100000111110111,
                                                                                        15'b101011111010100}};


key: 16, hash:13, tables: 32
localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,

                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = '{'{16'b1100001000100101,
                                                                                        16'b0001010001000101,
                                                                                        16'b1111101010111111,
                                                                                        16'b0011101010011001,
                                                                                        16'b1011001010100100,
                                                                                        16'b0010000100001101,
                                                                                        16'b0111011101010100,
                                                                                        16'b1001101011000000,
                                                                                        16'b0001101110111001,
                                                                                        16'b1001011101011010,
                                                                                        16'b0101111111100001,
                                                                                        16'b0101010111011110,
                                                                                        16'b0000000001101001},

                                                                                      '{16'b0111011100010010,
                                                                                        16'b0010001100100010,
                                                                                        16'b1011110011010100,
                                                                                        16'b1101001101011100,
                                                                                        16'b1010101001111110,
                                                                                        16'b0110111010111100,
                                                                                        16'b1011111001111001,
                                                                                        16'b0111000111111010,
                                                                                        16'b1111001001111100,
                                                                                        16'b0011001101100111,
                                                                                        16'b1101011101101111,
                                                                                        16'b1110000100000001,
                                                                                        16'b0111000001011001},

                                                                                      '{16'b1111100011000111,
                                                                                        16'b0110101011110010,
                                                                                        16'b1111100111000100,
                                                                                        16'b0001111001101100,
                                                                                        16'b1011100011011010,
                                                                                        16'b1111000010100000,
                                                                                        16'b1100100000111010,
                                                                                        16'b0100001000111000,
                                                                                        16'b1001001101101000,
                                                                                        16'b1100111011100000,
                                                                                        16'b1011010001010111,
                                                                                        16'b0101000101010001,
                                                                                        16'b1001101000000101}, 

                                                                                      '{16'b0001110100101110,
                                                                                        16'b1000000010100111,
                                                                                        16'b0010000100100011,
                                                                                        16'b0000110011011010,
                                                                                        16'b1001000001100011,
                                                                                        16'b1111011011101111,
                                                                                        16'b1001100111100110,
                                                                                        16'b1101010001000111,
                                                                                        16'b1111110011001101,
                                                                                        16'b1010000011111010,
                                                                                        16'b1110010110101001,
                                                                                        16'b0011111001000011,
                                                                                        16'b0101011100010100},

                                                                                      '{16'b1010001011010100,
                                                                                        16'b1101000100001100,
                                                                                        16'b0100000110110011,
                                                                                        16'b1010101001001010,
                                                                                        16'b0101101101001011,
                                                                                        16'b0011101000101001,
                                                                                        16'b1101011111010001,
                                                                                        16'b0100011001011100,
                                                                                        16'b1001001100100011,
                                                                                        16'b1111000101011110,
                                                                                        16'b1110100110011100,
                                                                                        16'b1001000001000001,
                                                                                        16'b1001000110010101},

                                                                                      '{16'b0000110011111001,
                                                                                        16'b0000000110100010,
                                                                                        16'b0100100000101010,
                                                                                        16'b0101111111110111,
                                                                                        16'b0101101110111010,
                                                                                        16'b0000010111010000,
                                                                                        16'b1001100011001011,
                                                                                        16'b0111000000101001,
                                                                                        16'b0001000001010110,
                                                                                        16'b1001001101101101,
                                                                                        16'b0100001001110000,
                                                                                        16'b0100101001000000,
                                                                                        16'b0011101111101111},

                                                                                      '{16'b0010101101100110,
                                                                                        16'b1110111010001110,
                                                                                        16'b0101111010101001,
                                                                                        16'b0010110110001101,
                                                                                        16'b0110100101011000,
                                                                                        16'b0011110111101111,
                                                                                        16'b0110111001111001,
                                                                                        16'b0010110011100100,
                                                                                        16'b0111110101110011,
                                                                                        16'b0111011011011001,
                                                                                        16'b0100011001101010,
                                                                                        16'b1000100111000001,
                                                                                        16'b0111001001010101},

                                                                                      '{16'b1000000010100001,
                                                                                        16'b0001100001101111,
                                                                                        16'b0011000000000100,
                                                                                        16'b0011110011111011,
                                                                                        16'b0000010100111001,
                                                                                        16'b0110001001101101,
                                                                                        16'b0011010011001011,
                                                                                        16'b1000110110100001,
                                                                                        16'b0100101001000100,
                                                                                        16'b0001010001010011,
                                                                                        16'b1000110101101000,
                                                                                        16'b0111100111110000,
                                                                                        16'b1110001011000110},

                                                                                      '{16'b1110010000111110,
                                                                                        16'b0110111001100100,
                                                                                        16'b1010111001010000,
                                                                                        16'b0100110000010110,
                                                                                        16'b1000000000001011,
                                                                                        16'b0111011000101001,
                                                                                        16'b1100000011101101,
                                                                                        16'b0110101001110111,
                                                                                        16'b1001001101100011,
                                                                                        16'b0100000111010101,
                                                                                        16'b0010110000010100,
                                                                                        16'b0110111000010101,
                                                                                        16'b0000110000101110},

                                                                                      '{16'b0110010110110001,
                                                                                        16'b1100010101100110,
                                                                                        16'b1101001010101101,
                                                                                        16'b1100000001100001,
                                                                                        16'b1100110011101101,
                                                                                        16'b1100101010000000,
                                                                                        16'b0100000011011010,
                                                                                        16'b0000010111010010,
                                                                                        16'b1011011110100100,
                                                                                        16'b1001011110010110,
                                                                                        16'b1101111001000010,
                                                                                        16'b0001101000001011,
                                                                                        16'b0000011011010011},

                                                                                      '{16'b0010111010001001,
                                                                                        16'b1010000110110100,
                                                                                        16'b1111110011000110,
                                                                                        16'b1000001101110101,
                                                                                        16'b1000110011111110,
                                                                                        16'b1111111001111000,
                                                                                        16'b0110010111001011,
                                                                                        16'b1001000010011101,
                                                                                        16'b0001000010000010,
                                                                                        16'b0100010011111111,
                                                                                        16'b0000001110100100,
                                                                                        16'b1110111110001101,
                                                                                        16'b0011100101011100},

                                                                                      '{16'b1001111011011111,
                                                                                        16'b0101111100101110,
                                                                                        16'b1111110000100000,
                                                                                        16'b1100000011000001,
                                                                                        16'b0100111100011111,
                                                                                        16'b0001100100100100,
                                                                                        16'b1111111111101000,
                                                                                        16'b1010000101011110,
                                                                                        16'b1111000010100010,
                                                                                        16'b0110100111010001,
                                                                                        16'b0111100010110111,
                                                                                        16'b1110001010010110,
                                                                                        16'b1000001100010000},

                                                                                      '{16'b0001000011001010,
                                                                                        16'b0100010000111001,
                                                                                        16'b0001011100111111,
                                                                                        16'b1100100100010001,
                                                                                        16'b1011100001001100,
                                                                                        16'b0100101110110101,
                                                                                        16'b0001001110001100,
                                                                                        16'b0000110101011110,
                                                                                        16'b1011110111110110,
                                                                                        16'b0010101110100100,
                                                                                        16'b0100100110001000,
                                                                                        16'b1000010001010000,
                                                                                        16'b1111000010001011},

                                                                                      '{16'b0101110111001110,
                                                                                        16'b0001110100100110,
                                                                                        16'b0010100110111011,
                                                                                        16'b1110001110101011,
                                                                                        16'b0011100001100110,
                                                                                        16'b1011010100110100,
                                                                                        16'b0010000001011111,
                                                                                        16'b0101000001101010,
                                                                                        16'b1100010101001000,
                                                                                        16'b1001111110100100,
                                                                                        16'b1101001111100001,
                                                                                        16'b1101010101110001,
                                                                                        16'b0000110010100101},

                                                                                      '{16'b1101110010101110,
                                                                                        16'b0000111010110001,
                                                                                        16'b1000100100110100,
                                                                                        16'b1111011110000100,
                                                                                        16'b1110111111011100,
                                                                                        16'b1101101000100111,
                                                                                        16'b0010001101110111,
                                                                                        16'b1111100101111101,
                                                                                        16'b0101101010010100,
                                                                                        16'b1011010111000100,
                                                                                        16'b1101111111010100,
                                                                                        16'b1010000111010101,
                                                                                        16'b0111001111010100},

                                                                                      '{16'b0000100001110001,
                                                                                        16'b0010110101111001,
                                                                                        16'b0001110101101110,
                                                                                        16'b1101001111101100,
                                                                                        16'b1101100001100000,
                                                                                        16'b0000010001011110,
                                                                                        16'b0010000011001001,
                                                                                        16'b0001011001110000,
                                                                                        16'b1111111101010000,
                                                                                        16'b1110101110101111,
                                                                                        16'b1110011011111111,
                                                                                        16'b1110001010010000,
                                                                                        16'b0101110111110001},

                                                                                      '{16'b1000010001000000,
                                                                                        16'b0010010001100111,
                                                                                        16'b1001001000101000,
                                                                                        16'b0111110000000111,
                                                                                        16'b1110110001001111,
                                                                                        16'b0110011010000001,
                                                                                        16'b1110100101010111,
                                                                                        16'b0111001000111011,
                                                                                        16'b1100010101011100,
                                                                                        16'b1011010011110110,
                                                                                        16'b1111111101110101,
                                                                                        16'b1000011100110110,
                                                                                        16'b0100000101010111},

                                                                                      '{16'b0001011011001001,
                                                                                        16'b0001011100110011,
                                                                                        16'b1111111101011010,
                                                                                        16'b1111000100011010,
                                                                                        16'b0011101010100101,
                                                                                        16'b1111000010110111,
                                                                                        16'b1011010010010101,
                                                                                        16'b1110111100100000,
                                                                                        16'b0011011110010101,
                                                                                        16'b0010111110110101,
                                                                                        16'b0001000000010010,
                                                                                        16'b0100000001110110,
                                                                                        16'b0100110010011000},

                                                                                      '{16'b1010110000101001,
                                                                                        16'b0001001010110010,
                                                                                        16'b1101010010101101,
                                                                                        16'b1110100110111001,
                                                                                        16'b0111111001110011,
                                                                                        16'b0100111000110100,
                                                                                        16'b1001101010011110,
                                                                                        16'b1100111011000011,
                                                                                        16'b1110111101100000,
                                                                                        16'b1011100001100100,
                                                                                        16'b0111000110101011,
                                                                                        16'b0101111101100001,
                                                                                        16'b1111101111100110},

                                                                                      '{16'b1110100000111011,
                                                                                        16'b1110011000011000,
                                                                                        16'b1001010011110000,
                                                                                        16'b1101110100101101,
                                                                                        16'b1010011100011010,
                                                                                        16'b0001101011000110,
                                                                                        16'b1011000101010001,
                                                                                        16'b0010100101010010,
                                                                                        16'b0010101001011100,
                                                                                        16'b1100011011110101,
                                                                                        16'b0010000100101000,
                                                                                        16'b0011100010000110,
                                                                                        16'b0010101011001111},

                                                                                      '{16'b1000100111000100,
                                                                                        16'b0111100000001110,
                                                                                        16'b0011010001010111,
                                                                                        16'b1100011010010011,
                                                                                        16'b0011101101100111,
                                                                                        16'b1110100011110001,
                                                                                        16'b0000010101101100,
                                                                                        16'b0000100000000111,
                                                                                        16'b1011111111100011,
                                                                                        16'b0111010101100011,
                                                                                        16'b0010101100111101,
                                                                                        16'b1111010011000000,
                                                                                        16'b0110001001110101},

                                                                                      '{16'b0011011110010101,
                                                                                        16'b0011010000001011,
                                                                                        16'b0010000100111111,
                                                                                        16'b0100111100010100,
                                                                                        16'b0111110110010010,
                                                                                        16'b0101110010001001,
                                                                                        16'b0011100111111001,
                                                                                        16'b1000000000001101,
                                                                                        16'b1011001100010100,
                                                                                        16'b0001101100010111,
                                                                                        16'b1011101001101111,
                                                                                        16'b1010100111100101,
                                                                                        16'b0111100111010110},

                                                                                      '{16'b1111000111101100,
                                                                                        16'b0100000100101000,
                                                                                        16'b1110000000001000,
                                                                                        16'b0110100000100111,
                                                                                        16'b0100000101011101,
                                                                                        16'b1011100000100010,
                                                                                        16'b1000101100110001,
                                                                                        16'b0000111011111010,
                                                                                        16'b0110011000100111,
                                                                                        16'b1000001011011111,
                                                                                        16'b1001001000010010,
                                                                                        16'b1101111100110101,
                                                                                        16'b1000101111011110},

                                                                                      '{16'b1101000000010011,
                                                                                        16'b0100100111010001,
                                                                                        16'b1000101001110111,
                                                                                        16'b1011110100010010,
                                                                                        16'b1011001010010010,
                                                                                        16'b1001101111011100,
                                                                                        16'b0100110011001011,
                                                                                        16'b0011110000101111,
                                                                                        16'b1000101101001000,
                                                                                        16'b0011000001101010,
                                                                                        16'b0001100100000101,
                                                                                        16'b0000110100010111,
                                                                                        16'b0000100000010010},

                                                                                      '{16'b0010100010000001,
                                                                                        16'b0011100111100100,
                                                                                        16'b1001100100001010,
                                                                                        16'b0011001000011001,
                                                                                        16'b0110000100110001,
                                                                                        16'b1110010111110111,
                                                                                        16'b1111011100110011,
                                                                                        16'b0000000001000111,
                                                                                        16'b0010110010101101,
                                                                                        16'b1111100011000111,
                                                                                        16'b1111101101110100,
                                                                                        16'b0010000000111110,
                                                                                        16'b1001001010000010},

                                                                                      '{16'b1101100100010000,
                                                                                        16'b0101111101011110,
                                                                                        16'b1000110111100010,
                                                                                        16'b0101111110001100,
                                                                                        16'b0011111011110000,
                                                                                        16'b0011111101110100,
                                                                                        16'b0011111011010001,
                                                                                        16'b1100011010000101,
                                                                                        16'b0001110011111100,
                                                                                        16'b1110101001111110,
                                                                                        16'b1101000100110110,
                                                                                        16'b0010111000111000,
                                                                                        16'b1101010100011011},

                                                                                      '{16'b1110111010011110,
                                                                                        16'b0100110001111000,
                                                                                        16'b1001010111100001,
                                                                                        16'b1000100011101000,
                                                                                        16'b0111101010001011,
                                                                                        16'b1000110000000000,
                                                                                        16'b0111000110101100,
                                                                                        16'b1101111110111101,
                                                                                        16'b0001011001100101,
                                                                                        16'b1010001001010111,
                                                                                        16'b1101011011101111,
                                                                                        16'b1100101101111111,
                                                                                        16'b1110010100100110},

                                                                                      '{16'b0101110010010101,
                                                                                        16'b1100100100000010,
                                                                                        16'b1000100100001111,
                                                                                        16'b0011000110010101,
                                                                                        16'b0001101100100111,
                                                                                        16'b0001001001010100,
                                                                                        16'b0001010000010101,
                                                                                        16'b1001100001001010,
                                                                                        16'b0010111000100101,
                                                                                        16'b0010110110100110,
                                                                                        16'b1100101100111011,
                                                                                        16'b1001011100001100,
                                                                                        16'b0110001101101010},

                                                                                      '{16'b0011100111100110,
                                                                                        16'b0011100101111011,
                                                                                        16'b0011010111100100,
                                                                                        16'b0001001001011011,
                                                                                        16'b1001110001000011,
                                                                                        16'b1100111101010010,
                                                                                        16'b0111100101000111,
                                                                                        16'b0000001101011000,
                                                                                        16'b1110011110111110,
                                                                                        16'b0010011111111001,
                                                                                        16'b0011010001010110,
                                                                                        16'b1111011000011110,
                                                                                        16'b1111000010000111},

                                                                                      '{16'b0001101111100001,
                                                                                        16'b0101010000000010,
                                                                                        16'b0110001001011100,
                                                                                        16'b0101010011100000,
                                                                                        16'b0100001010101100,
                                                                                        16'b0001011011111010,
                                                                                        16'b1000111010111101,
                                                                                        16'b0010100100101010,
                                                                                        16'b0001010101010101,
                                                                                        16'b0010110111100010,
                                                                                        16'b1010010111011101,
                                                                                        16'b1000000110011001,
                                                                                        16'b1110011011010010},
                                                                                    
                                                                                    
                                                                                    
                                                                                      '{16'b1000111010011100,
                                                                                        16'b1011011111101101,
                                                                                        16'b1100101100001111,
                                                                                        16'b1010111010000111,
                                                                                        16'b0011010111001000,
                                                                                        16'b0000100100011000,
                                                                                        16'b0100110100011100,
                                                                                        16'b1100000000000011,
                                                                                        16'b0110101100010110,
                                                                                        16'b1110111100101011,
                                                                                        16'b0011110011111110,
                                                                                        16'b1101100100101101,
                                                                                        16'b0010110101110011},

                                                                                      '{16'b1010101010011001,
                                                                                        16'b1010000001110001,
                                                                                        16'b0001110010000101,
                                                                                        16'b0110001111010001,
                                                                                        16'b1111011101000111,
                                                                                        16'b1100100011110111,
                                                                                        16'b0010010110011100,
                                                                                        16'b1011101010111110,
                                                                                        16'b1101101000001101,
                                                                                        16'b1000110000010111,
                                                                                        16'b0011010011110100,
                                                                                        16'b0111100100000110,
                                                                                        16'b1111110110000011}};









key: 16, hash:12, tables: 32
localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd12,32'd12,32'd12,32'd12,
                                                            32'd12,32'd12,32'd12,32'd12,
                                                            32'd12,32'd12,32'd12,32'd12,
                                                            32'd12,32'd12,32'd12,32'd12,

                                                            32'd12,32'd12,32'd12,32'd12,
                                                            32'd12,32'd12,32'd12,32'd12,
                                                            32'd12,32'd12,32'd12,32'd12,
                                                            32'd12,32'd12,32'd12,32'd12};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = '{'{16'b1100001000100101,
                                                                                      16'b0001010001000101,
                                                                                      16'b1111101010111111,
                                                                                      16'b0011101010011001,
                                                                                      16'b1011001010100100,
                                                                                      16'b0010000100001101,
                                                                                      16'b0111011101010100,
                                                                                      16'b1001101011000000,
                                                                                      16'b0001101110111001,
                                                                                      16'b1001011101011010,
                                                                                      16'b0101111111100001,
                                                                                      16'b0000000001101001},

                                                                                    '{16'b0111011100010010,
                                                                                      16'b0010001100100010,
                                                                                      16'b1011110011010100,
                                                                                      16'b1101001101011100,
                                                                                      16'b1010101001111110,
                                                                                      16'b0110111010111100,
                                                                                      16'b1011111001111001,
                                                                                      16'b0111000111111010,
                                                                                      16'b1111001001111100,
                                                                                      16'b0011001101100111,
                                                                                      16'b1101011101101111,
                                                                                      16'b0111000001011001},

                                                                                    '{16'b1111100011000111,
                                                                                      16'b0110101011110010,
                                                                                      16'b1111100111000100,
                                                                                      16'b0001111001101100,
                                                                                      16'b1011100011011010,
                                                                                      16'b1111000010100000,
                                                                                      16'b1100100000111010,
                                                                                      16'b0100001000111000,
                                                                                      16'b1001001101101000,
                                                                                      16'b1100111011100000,
                                                                                      16'b1011010001010111,
                                                                                      16'b1001101000000101}, 

                                                                                    '{16'b0001110100101110,
                                                                                      16'b1000000010100111,
                                                                                      16'b0010000100100011,
                                                                                      16'b0000110011011010,
                                                                                      16'b1001000001100011,
                                                                                      16'b1111011011101111,
                                                                                      16'b1001100111100110,
                                                                                      16'b1101010001000111,
                                                                                      16'b1111110011001101,
                                                                                      16'b1010000011111010,
                                                                                      16'b1110010110101001,
                                                                                      16'b0101011100010100},

                                                                                    '{16'b1010001011010100,
                                                                                      16'b1101000100001100,
                                                                                      16'b0100000110110011,
                                                                                      16'b1010101001001010,
                                                                                      16'b0101101101001011,
                                                                                      16'b0011101000101001,
                                                                                      16'b1101011111010001,
                                                                                      16'b0100011001011100,
                                                                                      16'b1001001100100011,
                                                                                      16'b1111000101011110,
                                                                                      16'b1110100110011100,
                                                                                      16'b1001000110010101},

                                                                                    '{16'b0000110011111001,
                                                                                      16'b0000000110100010,
                                                                                      16'b0100100000101010,
                                                                                      16'b0101111111110111,
                                                                                      16'b0101101110111010,
                                                                                      16'b0000010111010000,
                                                                                      16'b1001100011001011,
                                                                                      16'b0111000000101001,
                                                                                      16'b0001000001010110,
                                                                                      16'b1001001101101101,
                                                                                      16'b0100001001110000,
                                                                                      16'b0011101111101111},

                                                                                    '{16'b0010101101100110,
                                                                                      16'b1110111010001110,
                                                                                      16'b0101111010101001,
                                                                                      16'b0010110110001101,
                                                                                      16'b0110100101011000,
                                                                                      16'b0011110111101111,
                                                                                      16'b0110111001111001,
                                                                                      16'b0010110011100100,
                                                                                      16'b0111110101110011,
                                                                                      16'b0111011011011001,
                                                                                      16'b0100011001101010,
                                                                                      16'b0111001001010101},

                                                                                    '{16'b1000000010100001,
                                                                                      16'b0001100001101111,
                                                                                      16'b0011000000000100,
                                                                                      16'b0011110011111011,
                                                                                      16'b0000010100111001,
                                                                                      16'b0110001001101101,
                                                                                      16'b0011010011001011,
                                                                                      16'b1000110110100001,
                                                                                      16'b0100101001000100,
                                                                                      16'b0001010001010011,
                                                                                      16'b1000110101101000,
                                                                                      16'b1110001011000110},

                                                                                    '{16'b1110010000111110,
                                                                                      16'b0110111001100100,
                                                                                      16'b1010111001010000,
                                                                                      16'b0100110000010110,
                                                                                      16'b1000000000001011,
                                                                                      16'b0111011000101001,
                                                                                      16'b1100000011101101,
                                                                                      16'b0110101001110111,
                                                                                      16'b1001001101100011,
                                                                                      16'b0100000111010101,
                                                                                      16'b0010110000010100,
                                                                                      16'b0000110000101110},

                                                                                    '{16'b0110010110110001,
                                                                                      16'b1100010101100110,
                                                                                      16'b1101001010101101,
                                                                                      16'b1100000001100001,
                                                                                      16'b1100110011101101,
                                                                                      16'b1100101010000000,
                                                                                      16'b0100000011011010,
                                                                                      16'b0000010111010010,
                                                                                      16'b1011011110100100,
                                                                                      16'b1001011110010110,
                                                                                      16'b1101111001000010,
                                                                                      16'b0000011011010011},

                                                                                    '{16'b0010111010001001,
                                                                                      16'b1010000110110100,
                                                                                      16'b1111110011000110,
                                                                                      16'b1000001101110101,
                                                                                      16'b1000110011111110,
                                                                                      16'b1111111001111000,
                                                                                      16'b0110010111001011,
                                                                                      16'b1001000010011101,
                                                                                      16'b0001000010000010,
                                                                                      16'b0100010011111111,
                                                                                      16'b0000001110100100,
                                                                                      16'b0011100101011100},

                                                                                    '{16'b1001111011011111,
                                                                                      16'b0101111100101110,
                                                                                      16'b1111110000100000,
                                                                                      16'b1100000011000001,
                                                                                      16'b0100111100011111,
                                                                                      16'b0001100100100100,
                                                                                      16'b1111111111101000,
                                                                                      16'b1010000101011110,
                                                                                      16'b1111000010100010,
                                                                                      16'b0110100111010001,
                                                                                      16'b0111100010110111,
                                                                                      16'b1000001100010000},

                                                                                    '{16'b0001000011001010,
                                                                                      16'b0100010000111001,
                                                                                      16'b0001011100111111,
                                                                                      16'b1100100100010001,
                                                                                      16'b1011100001001100,
                                                                                      16'b0100101110110101,
                                                                                      16'b0001001110001100,
                                                                                      16'b0000110101011110,
                                                                                      16'b1011110111110110,
                                                                                      16'b0010101110100100,
                                                                                      16'b0100100110001000,
                                                                                      16'b1111000010001011},

                                                                                    '{16'b0101110111001110,
                                                                                      16'b0001110100100110,
                                                                                      16'b0010100110111011,
                                                                                      16'b1110001110101011,
                                                                                      16'b0011100001100110,
                                                                                      16'b1011010100110100,
                                                                                      16'b0010000001011111,
                                                                                      16'b0101000001101010,
                                                                                      16'b1100010101001000,
                                                                                      16'b1001111110100100,
                                                                                      16'b1101001111100001,
                                                                                      16'b0000110010100101},

                                                                                    '{16'b1101110010101110,
                                                                                      16'b0000111010110001,
                                                                                      16'b1000100100110100,
                                                                                      16'b1111011110000100,
                                                                                      16'b1110111111011100,
                                                                                      16'b1101101000100111,
                                                                                      16'b0010001101110111,
                                                                                      16'b1111100101111101,
                                                                                      16'b0101101010010100,
                                                                                      16'b1011010111000100,
                                                                                      16'b1101111111010100,
                                                                                      16'b0111001111010100},

                                                                                    '{16'b0000100001110001,
                                                                                      16'b0010110101111001,
                                                                                      16'b0001110101101110,
                                                                                      16'b1101001111101100,
                                                                                      16'b1101100001100000,
                                                                                      16'b0000010001011110,
                                                                                      16'b0010000011001001,
                                                                                      16'b0001011001110000,
                                                                                      16'b1111111101010000,
                                                                                      16'b1110101110101111,
                                                                                      16'b1110011011111111,
                                                                                      16'b0101110111110001},

                                                                                    '{16'b1000010001000000,
                                                                                      16'b0010010001100111,
                                                                                      16'b1001001000101000,
                                                                                      16'b0111110000000111,
                                                                                      16'b1110110001001111,
                                                                                      16'b0110011010000001,
                                                                                      16'b1110100101010111,
                                                                                      16'b0111001000111011,
                                                                                      16'b1100010101011100,
                                                                                      16'b1011010011110110,
                                                                                      16'b1111111101110101,
                                                                                      16'b0100000101010111},

                                                                                    '{16'b0001011011001001,
                                                                                      16'b0001011100110011,
                                                                                      16'b1111111101011010,
                                                                                      16'b1111000100011010,
                                                                                      16'b0011101010100101,
                                                                                      16'b1111000010110111,
                                                                                      16'b1011010010010101,
                                                                                      16'b1110111100100000,
                                                                                      16'b0011011110010101,
                                                                                      16'b0010111110110101,
                                                                                      16'b0001000000010010,
                                                                                      16'b0100110010011000},

                                                                                    '{16'b1010110000101001,
                                                                                      16'b0001001010110010,
                                                                                      16'b1101010010101101,
                                                                                      16'b1110100110111001,
                                                                                      16'b0111111001110011,
                                                                                      16'b0100111000110100,
                                                                                      16'b1001101010011110,
                                                                                      16'b1100111011000011,
                                                                                      16'b1110111101100000,
                                                                                      16'b1011100001100100,
                                                                                      16'b0111000110101011,
                                                                                      16'b1111101111100110},

                                                                                    '{16'b1110100000111011,
                                                                                      16'b1110011000011000,
                                                                                      16'b1001010011110000,
                                                                                      16'b1101110100101101,
                                                                                      16'b1010011100011010,
                                                                                      16'b0001101011000110,
                                                                                      16'b1011000101010001,
                                                                                      16'b0010100101010010,
                                                                                      16'b0010101001011100,
                                                                                      16'b1100011011110101,
                                                                                      16'b0010000100101000,
                                                                                      16'b0010101011001111},

                                                                                    '{16'b1000100111000100,
                                                                                      16'b0111100000001110,
                                                                                      16'b0011010001010111,
                                                                                      16'b1100011010010011,
                                                                                      16'b0011101101100111,
                                                                                      16'b1110100011110001,
                                                                                      16'b0000010101101100,
                                                                                      16'b0000100000000111,
                                                                                      16'b1011111111100011,
                                                                                      16'b0111010101100011,
                                                                                      16'b0010101100111101,
                                                                                      16'b0110001001110101},

                                                                                    '{16'b0011011110010101,
                                                                                      16'b0011010000001011,
                                                                                      16'b0010000100111111,
                                                                                      16'b0100111100010100,
                                                                                      16'b0111110110010010,
                                                                                      16'b0101110010001001,
                                                                                      16'b0011100111111001,
                                                                                      16'b1000000000001101,
                                                                                      16'b1011001100010100,
                                                                                      16'b0001101100010111,
                                                                                      16'b1011101001101111,
                                                                                      16'b0111100111010110},

                                                                                    '{16'b1111000111101100,
                                                                                      16'b0100000100101000,
                                                                                      16'b1110000000001000,
                                                                                      16'b0110100000100111,
                                                                                      16'b0100000101011101,
                                                                                      16'b1011100000100010,
                                                                                      16'b1000101100110001,
                                                                                      16'b0000111011111010,
                                                                                      16'b0110011000100111,
                                                                                      16'b1000001011011111,
                                                                                      16'b1001001000010010,
                                                                                      16'b1000101111011110},

                                                                                    '{16'b1101000000010011,
                                                                                      16'b0100100111010001,
                                                                                      16'b1000101001110111,
                                                                                      16'b1011110100010010,
                                                                                      16'b1011001010010010,
                                                                                      16'b1001101111011100,
                                                                                      16'b0100110011001011,
                                                                                      16'b0011110000101111,
                                                                                      16'b1000101101001000,
                                                                                      16'b0011000001101010,
                                                                                      16'b0001100100000101,
                                                                                      16'b0000100000010010},

                                                                                    '{16'b0010100010000001,
                                                                                      16'b0011100111100100,
                                                                                      16'b1001100100001010,
                                                                                      16'b0011001000011001,
                                                                                      16'b0110000100110001,
                                                                                      16'b1110010111110111,
                                                                                      16'b1111011100110011,
                                                                                      16'b0000000001000111,
                                                                                      16'b0010110010101101,
                                                                                      16'b1111100011000111,
                                                                                      16'b1111101101110100,
                                                                                      16'b1001001010000010},

                                                                                    '{16'b1101100100010000,
                                                                                      16'b0101111101011110,
                                                                                      16'b1000110111100010,
                                                                                      16'b0101111110001100,
                                                                                      16'b0011111011110000,
                                                                                      16'b0011111101110100,
                                                                                      16'b0011111011010001,
                                                                                      16'b1100011010000101,
                                                                                      16'b0001110011111100,
                                                                                      16'b1110101001111110,
                                                                                      16'b1101000100110110,
                                                                                      16'b1101010100011011},

                                                                                    '{16'b1110111010011110,
                                                                                      16'b0100110001111000,
                                                                                      16'b1001010111100001,
                                                                                      16'b1000100011101000,
                                                                                      16'b0111101010001011,
                                                                                      16'b1000110000000000,
                                                                                      16'b0111000110101100,
                                                                                      16'b1101111110111101,
                                                                                      16'b0001011001100101,
                                                                                      16'b1010001001010111,
                                                                                      16'b1101011011101111,
                                                                                      16'b1110010100100110},

                                                                                    '{16'b0101110010010101,
                                                                                      16'b1100100100000010,
                                                                                      16'b1000100100001111,
                                                                                      16'b0011000110010101,
                                                                                      16'b0001101100100111,
                                                                                      16'b0001001001010100,
                                                                                      16'b0001010000010101,
                                                                                      16'b1001100001001010,
                                                                                      16'b0010111000100101,
                                                                                      16'b0010110110100110,
                                                                                      16'b1100101100111011,
                                                                                      16'b0110001101101010},

                                                                                    '{16'b0011100111100110,
                                                                                      16'b0011100101111011,
                                                                                      16'b0011010111100100,
                                                                                      16'b0001001001011011,
                                                                                      16'b1001110001000011,
                                                                                      16'b1100111101010010,
                                                                                      16'b0111100101000111,
                                                                                      16'b0000001101011000,
                                                                                      16'b1110011110111110,
                                                                                      16'b0010011111111001,
                                                                                      16'b0011010001010110,
                                                                                      16'b1111000010000111},

                                                                                    '{16'b0001101111100001,
                                                                                      16'b0101010000000010,
                                                                                      16'b0110001001011100,
                                                                                      16'b0101010011100000,
                                                                                      16'b0100001010101100,
                                                                                      16'b0001011011111010,
                                                                                      16'b1000111010111101,
                                                                                      16'b0010100100101010,
                                                                                      16'b0001010101010101,
                                                                                      16'b0010110111100010,
                                                                                      16'b1010010111011101,
                                                                                      16'b1110011011010010},
                                                                                  
                                                                                  
                                                                                  
                                                                                    '{16'b1000111010011100,
                                                                                      16'b1011011111101101,
                                                                                      16'b1100101100001111,
                                                                                      16'b1010111010000111,
                                                                                      16'b0011010111001000,
                                                                                      16'b0000100100011000,
                                                                                      16'b0100110100011100,
                                                                                      16'b1100000000000011,
                                                                                      16'b0110101100010110,
                                                                                      16'b1110111100101011,
                                                                                      16'b0011110011111110,
                                                                                      16'b0010110101110011},

                                                                                    '{16'b1010101010011001,
                                                                                      16'b1010000001110001,
                                                                                      16'b0001110010000101,
                                                                                      16'b0110001111010001,
                                                                                      16'b1111011101000111,
                                                                                      16'b1100100011110111,
                                                                                      16'b0010010110011100,
                                                                                      16'b1011101010111110,
                                                                                      16'b1101101000001101,
                                                                                      16'b1000110000010111,
                                                                                      16'b0011010011110100,
                                                                                      16'b1111110110000011}};







key: 16, hash:14, tables: 8
localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd14,32'd14,32'd14,32'd14,
                                                             32'd14,32'd14,32'd14,32'd14};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = 
                                                                                    '{'{16'b1100001000100101,
                                                                                        16'b0001010001000101,
                                                                                        16'b1111101010111111,
                                                                                        16'b0011101010011001,
                                                                                        16'b1011001010100100,
                                                                                        16'b0010000100001101,
                                                                                        16'b0111011101010100,
                                                                                        16'b0100000111101111,
                                                                                        16'b0010010101000011,
                                                                                        16'b1001101011000000,
                                                                                        16'b0001101110111001,
                                                                                        16'b1001011101011010,
                                                                                        16'b0101111111100001,
                                                                                        16'b0000000001101001},
                           
                                                                                      '{16'b0111011100010010,
                                                                                        16'b0010001100100010,
                                                                                        16'b1011110011010100,
                                                                                        16'b1101111000001000,
                                                                                        16'b0110101001001000,
                                                                                        16'b1101001101011100,
                                                                                        16'b1010101001111110,
                                                                                        16'b0110111010111100,
                                                                                        16'b1011111001111001,
                                                                                        16'b0111000111111010,
                                                                                        16'b1111001001111100,
                                                                                        16'b0011001101100111,
                                                                                        16'b1101011101101111,
                                                                                        16'b0111000001011001},
                           
                                                                                      '{16'b1111100011000111,
                                                                                        16'b0110101011110010,
                                                                                        16'b1111100111000100,
                                                                                        16'b0001111001101100,
                                                                                        16'b0011000001101001,
                                                                                        16'b1010001110111010,
                                                                                        16'b1011100011011010,
                                                                                        16'b1111000010100000,
                                                                                        16'b1100100000111010,
                                                                                        16'b0100001000111000,
                                                                                        16'b1001001101101000,
                                                                                        16'b1100111011100000,
                                                                                        16'b1011010001010111,
                                                                                        16'b1001101000000101}, 
                           
                                                                                      '{16'b0001110100101110,
                                                                                        16'b1000000010100111,
                                                                                        16'b0010000100100011,
                                                                                        16'b0000110011011010,
                                                                                        16'b0100011111000111,
                                                                                        16'b0011110010010100,
                                                                                        16'b1001000001100011,
                                                                                        16'b1111011011101111,
                                                                                        16'b1001100111100110,
                                                                                        16'b1101010001000111,
                                                                                        16'b1111110011001101,
                                                                                        16'b1010000011111010,
                                                                                        16'b1110010110101001,
                                                                                        16'b0101011100010100},
                           
                                                                                      '{16'b1010001011010100,
                                                                                        16'b1101000100001100,
                                                                                        16'b0100000110110011,
                                                                                        16'b1010101001001010,
                                                                                        16'b0101101101001011,
                                                                                        16'b0011101000101001,
                                                                                        16'b1101011111010001,
                                                                                        16'b0101000100100011,
                                                                                        16'b0111010011111010,
                                                                                        16'b0100011001011100,
                                                                                        16'b1001001100100011,
                                                                                        16'b1111000101011110,
                                                                                        16'b1110100110011100,
                                                                                        16'b1001000110010101},
                           
                                                                                      '{16'b0000110011111001,
                                                                                        16'b0000000110100010,
                                                                                        16'b0100100000101010,
                                                                                        16'b0101111111110111,
                                                                                        16'b0101101110111010,
                                                                                        16'b1110000010000100,
                                                                                        16'b1100110111011110,
                                                                                        16'b0000010111010000,
                                                                                        16'b1001100011001011,
                                                                                        16'b0111000000101001,
                                                                                        16'b0001000001010110,
                                                                                        16'b1001001101101101,
                                                                                        16'b0100001001110000,
                                                                                        16'b0011101111101111},
                           
                                                                                      '{16'b0010101101100110,
                                                                                        16'b1110111010001110,
                                                                                        16'b0101111010101001,
                                                                                        16'b0010110110001101,
                                                                                        16'b0110100101011000,
                                                                                        16'b1001101100101100,
                                                                                        16'b0101111001001101,
                                                                                        16'b0011110111101111,
                                                                                        16'b0110111001111001,
                                                                                        16'b0010110011100100,
                                                                                        16'b0111110101110011,
                                                                                        16'b0111011011011001,
                                                                                        16'b0100011001101010,
                                                                                        16'b0111001001010101},
                           
                                                                                      '{16'b1000000010100001,
                                                                                        16'b0001100001101111,
                                                                                        16'b0011000000000100,
                                                                                        16'b0011110011111011,
                                                                                        16'b1001111100111000,
                                                                                        16'b0101001100100010,
                                                                                        16'b0000010100111001,
                                                                                        16'b0110001001101101,
                                                                                        16'b0011010011001011,
                                                                                        16'b1000110110100001,
                                                                                        16'b0100101001000100,
                                                                                        16'b0001010001010011,
                                                                                        16'b1000110101101000,
                                                                                        16'b1110001011000110}};






key: 16, hash:13, tables: 16
localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13,
                                                             32'd13,32'd13,32'd13,32'd13};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = 
                                                         '{'{16'b1000010001000000,
                                                             16'b0010010001100111,
                                                             16'b1001001000101000,
                                                             16'b0111110000000111,
                                                             16'b1110110001001111,
                                                             16'b0110011010000001,
                                                             16'b1110100101010111,
                                                             16'b0111001000111011,
                                                             16'b1100010101011100,
                                                             16'b1011010011110110,
                                                             16'b1111111101110101,
                                                             16'b0110111100010100,
                                                             16'b0100000101010111},

                                                           '{16'b0001011011001001,
                                                             16'b0001011100110011,
                                                             16'b1111111101011010,
                                                             16'b1111000100011010,
                                                             16'b0011101010100101,
                                                             16'b1111000010110111,
                                                             16'b1011010010010101,
                                                             16'b1110111100100000,
                                                             16'b0011011110010101,
                                                             16'b0010111110110101,
                                                             16'b0001000000010010,
                                                             16'b0110010111100000,
                                                             16'b0100110010011000},

                                                           '{16'b1010110000101001,
                                                             16'b0001001010110010,
                                                             16'b1101010010101101,
                                                             16'b1110100110111001,
                                                             16'b0111111001110011,
                                                             16'b0100111000110100,
                                                             16'b1001101010011110,
                                                             16'b1100111011000011,
                                                             16'b1110111101100000,
                                                             16'b1011100001100100,
                                                             16'b0111000110101011,
                                                             16'b0101011010000100,
                                                             16'b1111101111100110},

                                                           '{16'b1110100000111011,
                                                             16'b1110011000011000,
                                                             16'b1001010011110000,
                                                             16'b1101110100101101,
                                                             16'b1010011100011010,
                                                             16'b0001101011000110,
                                                             16'b1011000101010001,
                                                             16'b0010100101010010,
                                                             16'b0010101001011100,
                                                             16'b1100011011110101,
                                                             16'b0010000100101000,
                                                             16'b1001000111000001,
                                                             16'b0010101011001111},

                                                           '{16'b1000100111000100,
                                                             16'b0111100000001110,
                                                             16'b0011010001010111,
                                                             16'b1100011010010011,
                                                             16'b0011101101100111,
                                                             16'b1110100011110001,
                                                             16'b0000010101101100,
                                                             16'b0000100000000111,
                                                             16'b1011111111100011,
                                                             16'b0111010101100011,
                                                             16'b0010101100111101,
                                                             16'b0100101111010011,
                                                             16'b0110001001110101},

                                                           '{16'b0011011110010101,
                                                             16'b0011010000001011,
                                                             16'b0010000100111111,
                                                             16'b0100111100010100,
                                                             16'b0111110110010010,
                                                             16'b0101110010001001,
                                                             16'b0011100111111001,
                                                             16'b1000000000001101,
                                                             16'b1011001100010100,
                                                             16'b0001101100010111,
                                                             16'b1011101001101111,
                                                             16'b1101011111010010,
                                                             16'b0111100111010110},

                                                           '{16'b1111000111101100,
                                                             16'b0100000100101000,
                                                             16'b1110000000001000,
                                                             16'b0110100000100111,
                                                             16'b0100000101011101,
                                                             16'b1011100000100010,
                                                             16'b1000101100110001,
                                                             16'b0000111011111010,
                                                             16'b0110011000100111,
                                                             16'b1000001011011111,
                                                             16'b1001001000010010,
                                                             16'b1110011000001011,
                                                             16'b1000101111011110},

                                                           '{16'b1101000000010011,
                                                             16'b0100100111010001,
                                                             16'b1000101001110111,
                                                             16'b1011110100010010,
                                                             16'b1011001010010010,
                                                             16'b1001101111011100,
                                                             16'b0100110011001011,
                                                             16'b0011110000101111,
                                                             16'b1000101101001000,
                                                             16'b0011000001101010,
                                                             16'b0001100100000101,
                                                             16'b1011111100100001,
                                                             16'b0000100000010010},

                                                           '{16'b0010100010000001,
                                                             16'b0011100111100100,
                                                             16'b1001100100001010,
                                                             16'b0011001000011001,
                                                             16'b0110000100110001,
                                                             16'b1110010111110111,
                                                             16'b1111011100110011,
                                                             16'b0000000001000111,
                                                             16'b0010110010101101,
                                                             16'b1111100011000111,
                                                             16'b1111101101110100,
                                                             16'b1111000111010001,
                                                             16'b1001001010000010},

                                                           '{16'b1101100100010000,
                                                             16'b0101111101011110,
                                                             16'b1000110111100010,
                                                             16'b0101111110001100,
                                                             16'b0011111011110000,
                                                             16'b0011111101110100,
                                                             16'b0011111011010001,
                                                             16'b1100011010000101,
                                                             16'b0001110011111100,
                                                             16'b1110101001111110,
                                                             16'b1101000100110110,
                                                             16'b1111000000001111,
                                                             16'b1101010100011011},

                                                           '{16'b1110111010011110,
                                                             16'b0100110001111000,
                                                             16'b1001010111100001,
                                                             16'b1000100011101000,
                                                             16'b0111101010001011,
                                                             16'b1000110000000000,
                                                             16'b0111000110101100,
                                                             16'b1101111110111101,
                                                             16'b0001011001100101,
                                                             16'b1010001001010111,
                                                             16'b1101011011101111,
                                                             16'b0101110010011110,
                                                             16'b1110010100100110},

                                                           '{16'b0101110010010101,
                                                             16'b1100100100000010,
                                                             16'b1000100100001111,
                                                             16'b0011000110010101,
                                                             16'b0001101100100111,
                                                             16'b0001001001010100,
                                                             16'b0001010000010101,
                                                             16'b1001100001001010,
                                                             16'b0010111000100101,
                                                             16'b0010110110100110,
                                                             16'b1100101100111011,
                                                             16'b0010100100100001,
                                                             16'b0110001101101010},

                                                           '{16'b0011100111100110,
                                                             16'b0011100101111011,
                                                             16'b0011010111100100,
                                                             16'b0001001001011011,
                                                             16'b1001110001000011,
                                                             16'b1100111101010010,
                                                             16'b0111100101000111,
                                                             16'b0000001101011000,
                                                             16'b1110011110111110,
                                                             16'b0010011111111001,
                                                             16'b0011010001010110,
                                                             16'b0000111100011000,
                                                             16'b1111000010000111},

                                                           '{16'b0001101111100001,
                                                             16'b0101010000000010,
                                                             16'b0110001001011100,
                                                             16'b0101010011100000,
                                                             16'b0100001010101100,
                                                             16'b0001011011111010,
                                                             16'b1000111010111101,
                                                             16'b0010100100101010,
                                                             16'b0001010101010101,
                                                             16'b0010110111100010,
                                                             16'b1010010111011101,
                                                             16'b1011110010111110,
                                                             16'b1110011011010010},
                                                         
                                                         
                                                         
                                                           '{16'b1000111010011100,
                                                             16'b1011011111101101,
                                                             16'b1100101100001111,
                                                             16'b1010111010000111,
                                                             16'b0011010111001000,
                                                             16'b0000100100011000,
                                                             16'b0100110100011100,
                                                             16'b1100000000000011,
                                                             16'b0110101100010110,
                                                             16'b1110111100101011,
                                                             16'b0011110011111110,
                                                             16'b1011110010111110,
                                                             16'b0010110101110011},

                                                           '{16'b1010101010011001,
                                                             16'b1010000001110001,
                                                             16'b0001110010000101,
                                                             16'b0110001111010001,
                                                             16'b1111011101000111,
                                                             16'b1100100011110111,
                                                             16'b0010010110011100,
                                                             16'b1011101010111110,
                                                             16'b1101101000001101,
                                                             16'b1000110000010111,
                                                             16'b0011010011110100,
                                                             16'b0101110101011001,
                                                             16'b1111110110000011}};