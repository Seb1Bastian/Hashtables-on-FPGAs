module matrix_generator #(parameter NUMBER_OF_TABLES = 4,
                          parameter HASH_ADR_WIDTH   = 5,
                          parameter KEY_WIDTH = 6)(
    output  wire  [NUMBER_OF_TABLES*HASH_ADR_WIDTH*KEY_WIDTH-1:0]  matrixes_o
); 

wire[KEY_WIDTH-1:0] logic_matrix[NUMBER_OF_TABLES-1:0][HASH_ADR_WIDTH-1:0];

localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd11,32'd11,32'd11,32'd11,
                                                             32'd11,32'd11,32'd11,32'd11};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = 
                                                                                    '{'{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001}, 
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001},
                           
                                                                                      '{32'b00000000000000000000010000000000,
                                                                                        32'b00000000000000000000001000000000,
                                                                                        32'b00000000000000000000000100000000,
                                                                                        32'b00000000000000000000000010000000,
                                                                                        32'b00000000000000000000000001000000,
                                                                                        32'b00000000000000000000000000100000,
                                                                                        32'b00000000000000000000000000010000,
                                                                                        32'b00000000000000000000000000001000,
                                                                                        32'b00000000000000000000000000000100,
                                                                                        32'b00000000000000000000000000000010,
                                                                                        32'b00000000000000000000000000000001}};
genvar i,j,l;
generate
    for (i = 0; i < NUMBER_OF_TABLES; i++) begin
        for (j = 0; j < HASH_ADR_WIDTH; j++) begin
            for (l = 0; l < KEY_WIDTH; l++) begin
                assign logic_matrix[i][j][l] = Q_MATRIX[i][j][l];
            end
        end
    end
endgenerate

generate
    for (i = 0; i < NUMBER_OF_TABLES; i++) begin
        for (j = 0; j < HASH_ADR_WIDTH; j++) begin
            assign matrixes_o[(i * HASH_ADR_WIDTH * KEY_WIDTH) + (j * KEY_WIDTH) +: KEY_WIDTH] = logic_matrix[i][j];
        end
    end
endgenerate

endmodule