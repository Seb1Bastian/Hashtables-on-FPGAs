key: 15, hash:10, tables: 10
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = '{'{15'b001001100011100,
                                                                                        15'b000000000100001,
                                                                                        15'b000000100011101,
                                                                                        15'b100010111010001,
                                                                                        15'b010000011110100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100010011000,
                                                                                        15'b100011100100110,
                                                                                        15'b011001000101000,
                                                                                        15'b111110001001010},
                                                                                    '{15'b010001011001001,
                                                                                        15'b001000000100000,
                                                                                        15'b001000010100101,
                                                                                        15'b011100010001000,
                                                                                        15'b100011110001111,
                                                                                        15'b001000101000100,
                                                                                        15'b000000000011000,
                                                                                        15'b011111000010000,
                                                                                        15'b000001000100101,
                                                                                        15'b000110000101101}, 
                                                                                    '{15'b000110100000110,
                                                                                        15'b101100110000100,
                                                                                        15'b010001001000111,
                                                                                        15'b001110010010100,
                                                                                        15'b101010010000100,
                                                                                        15'b000101101011001,
                                                                                        15'b001011000010010,
                                                                                        15'b110010100010010,
                                                                                        15'b001000100010110,
                                                                                        15'b110001100010000},

                                                                                    '{15'b001001000011100,
                                                                                        15'b101100000100001,
                                                                                        15'b011000001011101,
                                                                                        15'b010010101010001,
                                                                                        15'b010110011010100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100011011000,
                                                                                        15'b100010001101110,
                                                                                        15'b111001000101000,
                                                                                        15'b110010101011010},
                                                                                    '{15'b010001011001011,
                                                                                        15'b001000000111000,
                                                                                        15'b001000010000101,
                                                                                        15'b011100010101000,
                                                                                        15'b111000110001111,
                                                                                        15'b001001001000100,
                                                                                        15'b010001100011000,
                                                                                        15'b011011000000111,
                                                                                        15'b011001010000110,
                                                                                        15'b100100110111001}, 
                                                                                    '{15'b011001100111110,
                                                                                        15'b110110100011010,
                                                                                        15'b001010101000000,
                                                                                        15'b100001101011100,
                                                                                        15'b011111111001000,
                                                                                        15'b110011101110101,
                                                                                        15'b101010110001001,
                                                                                        15'b010000010111011,
                                                                                        15'b000110100110010,
                                                                                        15'b100101011011101},
                                                                                    '{15'b101010001011100,
                                                                                        15'b010110101101000,
                                                                                        15'b111010010000101,
                                                                                        15'b110000111111011,
                                                                                        15'b101100110111000,
                                                                                        15'b110001001010111,
                                                                                        15'b101100110000001,
                                                                                        15'b101001110110010,
                                                                                        15'b010101010111100,
                                                                                        15'b000101011011010},
                                                                                    '{15'b011001000000100,
                                                                                        15'b101100001010000,
                                                                                        15'b000000110101100,
                                                                                        15'b101111110100100,
                                                                                        15'b010011100111000,
                                                                                        15'b001100000001010,
                                                                                        15'b000111101110110,
                                                                                        15'b101010010001011,
                                                                                        15'b000101010110101,
                                                                                        15'b001100011001111}, 
                                                                                    '{15'b110111111011111,
                                                                                        15'b100100111110001,
                                                                                        15'b001011111110100,
                                                                                        15'b110100001010110,
                                                                                        15'b010110011110010,
                                                                                        15'b010001001110100,
                                                                                        15'b100110001011101,
                                                                                        15'b010111111111001,
                                                                                        15'b101000001100001,
                                                                                        15'b110011010111010},
                                                                                    '{15'b101010100101001,
                                                                                        15'b101011111101011,
                                                                                        15'b000011011010100,
                                                                                        15'b110011000101011,
                                                                                        15'b111011000111011,
                                                                                        15'b000001101000100,
                                                                                        15'b111000011100000,
                                                                                        15'b110011010010111,
                                                                                        15'b100000111110111,
                                                                                        15'b101011111010100}};


key: 15, hash:13, tables: 10
localparam integer HASH_TABLE_SIZE[NUMBER_OF_TABLES-1:0] = '{32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13,32'd13};
localparam [KEY_WIDTH-1:0] Q_MATRIX[NUMBER_OF_TABLES-1:0][HASH_TABLE_SIZE[0]-1:0] = '{'{15'b001001100011100,
                                                                                        15'b000000000100001,
                                                                                        15'b000000100011101,
                                                                                        15'b100010111010001,
                                                                                        15'b010000011110100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100010011000,
                                                                                        15'b010011101111010,
                                                                                        15'b100001111000101,
                                                                                        15'b101101111001001,
                                                                                        15'b100011100100110,
                                                                                        15'b011001000101000,
                                                                                        15'b111110001001010},
                                                                                    '{15'b010001011001001,
                                                                                        15'b001000000100000,
                                                                                        15'b001000010100101,
                                                                                        15'b011100010001000,
                                                                                        15'b011100000101100,
                                                                                        15'b001001110100101,
                                                                                        15'b101010010001000,
                                                                                        15'b100011110001111,
                                                                                        15'b001000101000100,
                                                                                        15'b000000000011000,
                                                                                        15'b011111000010000,
                                                                                        15'b000001000100101,
                                                                                        15'b000110000101101}, 
                                                                                    '{15'b000110100000110,
                                                                                        15'b101100110000100,
                                                                                        15'b010001001000111,
                                                                                        15'b001110010010100,
                                                                                        15'b101010010000100,
                                                                                        15'b000101101011001,
                                                                                        15'b001011000010010,
                                                                                        15'b110010100010010,
                                                                                        15'b001000100010110,
                                                                                        15'b001011001110010,
                                                                                        15'b110110101110010,
                                                                                        15'b001011100000110,
                                                                                        15'b110001100010000},

                                                                                    '{15'b001001000011100,
                                                                                        15'b101100000100001,
                                                                                        15'b011000001011101,
                                                                                        15'b010010101010001,
                                                                                        15'b101111000100001,
                                                                                        15'b011001101011101,
                                                                                        15'b110010101010001,
                                                                                        15'b010110011010100,
                                                                                        15'b100011001000101,
                                                                                        15'b101100011011000,
                                                                                        15'b100010001101110,
                                                                                        15'b111001000101000,
                                                                                        15'b110010101011010},
                                                                                    '{15'b010001011001011,
                                                                                        15'b001000000111000,
                                                                                        15'b001000010000101,
                                                                                        15'b011100010101000,
                                                                                        15'b111000111001111,
                                                                                        15'b010110110101000,
                                                                                        15'b111000111010111,
                                                                                        15'b001001001000100,
                                                                                        15'b001001001000100,
                                                                                        15'b010001100011000,
                                                                                        15'b011011000000111,
                                                                                        15'b011001010000110,
                                                                                        15'b100100110111001}, 
                                                                                    '{15'b011001100111110,
                                                                                        15'b110110100011010,
                                                                                        15'b001010101000000,
                                                                                        15'b100001101011100,
                                                                                        15'b011111111001000,
                                                                                        15'b110011101110101,
                                                                                        15'b101010110001001,
                                                                                        15'b101011101110101,
                                                                                        15'b101010110110001,
                                                                                        15'b010011010110011,
                                                                                        15'b010000010111011,
                                                                                        15'b000110100110010,
                                                                                        15'b100101011011101},
                                                                                    '{15'b101010001011100,
                                                                                        15'b010110101101000,
                                                                                        15'b101101110101001,
                                                                                        15'b110101001010110,
                                                                                        15'b101000110011011,
                                                                                        15'b111010010000101,
                                                                                        15'b110000111111011,
                                                                                        15'b101100110111000,
                                                                                        15'b110001001010111,
                                                                                        15'b101100110000001,
                                                                                        15'b101001110110010,
                                                                                        15'b010101010111100,
                                                                                        15'b000101011011010},
                                                                                    '{15'b011001000000100,
                                                                                        15'b101100001010000,
                                                                                        15'b000000110101100,
                                                                                        15'b101111110100100,
                                                                                        15'b010011100111000,
                                                                                        15'b110011110110001,
                                                                                        15'b101101010001010,
                                                                                        15'b100110101110110,
                                                                                        15'b001100000001010,
                                                                                        15'b000111101110110,
                                                                                        15'b101010010001011,
                                                                                        15'b000101010110101,
                                                                                        15'b001100011001111}, 
                                                                                    '{15'b110111111011111,
                                                                                        15'b100100111110001,
                                                                                        15'b110110010110010,
                                                                                        15'b011001001100101,
                                                                                        15'b100101001011101,
                                                                                        15'b001011111110100,
                                                                                        15'b110100001010110,
                                                                                        15'b010110011110010,
                                                                                        15'b010001001110100,
                                                                                        15'b100110001011101,
                                                                                        15'b010111111111001,
                                                                                        15'b101000001100001,
                                                                                        15'b110011010111010},
                                                                                    '{15'b101010100101001,
                                                                                        15'b101011111101011,
                                                                                        15'b000011011010100,
                                                                                        15'b110011000101011,
                                                                                        15'b111011000111011,
                                                                                        15'b101011011100000,
                                                                                        15'b110111010010111,
                                                                                        15'b100100100110111,
                                                                                        15'b000001101000100,
                                                                                        15'b111000011100000,
                                                                                        15'b110011010010111,
                                                                                        15'b100000111110111,
                                                                                        15'b101011111010100}};